module dram
(
  input i_clk, 
  input i_rst,
  input i_wr_en,
  input [31:0] i_wr_addr,
  input [31:0] i_wr_data, 
  input i_rd_en,   
  input [31:0] i_rd_addr, 

  output reg [31:0] o_rd_data,
  output reg o_valid
);


// Here for the fake memory, only 4 will be implemented
reg [31:0] REG [0:9999];


always @ (posedge i_clk or negedge i_rst) begin
	if (~i_rst) begin
		o_rd_data <= 0;
	  	o_valid <= 0;
	end
	else begin
	  if(i_rd_en) begin 
	  	// if (i_rd_addr<16'd6145) o_rd_data <= REG[i_rd_addr];
	  	// else begin
	  	// 	o_rd_data <= i_rd_addr[31:0];
	  	// end
	  	o_rd_data <= {REG[i_rd_addr][7:0],REG[i_rd_addr][15:8],REG[i_rd_addr][23:16],REG[i_rd_addr][31:24]};
	  	// o_rd_data <= {16'b0,i_rd_addr};
	  	o_valid <= 1;
	  end
	  else begin 
	  	o_rd_data <= 32'bx;
	  	o_valid <= 0;
	  end
	end
end


always @ (posedge i_clk or negedge i_rst) begin
	if (~i_rst) begin
////////////////////////////////////////////////////
//// IFMAP
////////////////////////////////////////////////////
REG[0] <= 32'b00000000000000000000000000000000;
REG[1] <= 32'b00000000000000000000000000000000;
REG[2] <= 32'b00000000000000000000000000000000;
REG[3] <= 32'b00000000000000000000000000000000;
REG[4] <= 32'b00000000000000100000000000000000;
REG[5] <= 32'b00000000000000000000000000000000;
REG[6] <= 32'b00000000000000000000000000000000;
REG[7] <= 32'b00000000000000000000000000000000;
REG[8] <= 32'b00000000000000000000010100000000;
REG[9] <= 32'b00000000000000000000000000000000;
REG[10] <= 32'b00000000000000000000000000000000;
REG[11] <= 32'b00000000000000000000010100000000;
REG[12] <= 32'b00000000000000000000000000000000;
REG[13] <= 32'b00000000000000000000000000000000;
REG[14] <= 32'b00000000000000000000000000000000;
REG[15] <= 32'b00000000000011000000000000000100;
REG[16] <= 32'b00000000000000000011111000101101;
REG[17] <= 32'b00000000000000000000000000000000;
REG[18] <= 32'b00000001000000000000000000000000;
REG[19] <= 32'b00010101000000000000011000110001;
REG[20] <= 32'b00000000000000000000000000000000;
REG[21] <= 32'b00001010000000000000000000000000;
REG[22] <= 32'b00000110000000000000000000001111;
REG[23] <= 32'b00010010000000000000000000000000;
REG[24] <= 32'b00000000000000000000000000000000;
REG[25] <= 32'b00000000000000000000000000000000;
REG[26] <= 32'b00000000000000000000000000000000;
REG[27] <= 32'b00000000000000000000000000000000;
REG[28] <= 32'b00000000000000000000000000000000;
REG[29] <= 32'b00100010000000000000010000010110;
REG[30] <= 32'b00000000000001000000000000000000;
REG[31] <= 32'b00000000000000000000000000000000;
REG[32] <= 32'b00000000000000000001101100000000;
REG[33] <= 32'b00000000010000110010100100000000;
REG[34] <= 32'b00000000000000000000000000001001;
REG[35] <= 32'b00000000000000000000001000000000;
REG[36] <= 32'b00000000000000000000000000000000;
REG[37] <= 32'b00000000000000000000000000000000;
REG[38] <= 32'b00000000000000000000000000000000;
REG[39] <= 32'b00000000000000000000000000000000;
REG[40] <= 32'b00000000000000000010000000000000;
REG[41] <= 32'b00000000000000100000000000000000;
REG[42] <= 32'b00000000000000000000000000000000;
REG[43] <= 32'b00000000000000000000000000000000;
REG[44] <= 32'b00000000000000000000011100000000;
REG[45] <= 32'b00010101000000000000000000000000;
REG[46] <= 32'b00000000000000000000000000000000;
REG[47] <= 32'b00000000000000000000000000000100;
REG[48] <= 32'b00000000000000000000000000000000;
REG[49] <= 32'b00000000000000000000000000000000;
REG[50] <= 32'b00000000000000000000000000000000;
REG[51] <= 32'b00000000000000000000000000000000;
REG[52] <= 32'b00010100000000000000000000000000;
REG[53] <= 32'b00010111000000000000000000000000;
REG[54] <= 32'b00000000000000000000000000000000;
REG[55] <= 32'b00001011000000110000000000000000;
REG[56] <= 32'b00000100000000000000000000000000;
REG[57] <= 32'b00000000000000000000000000000000;
REG[58] <= 32'b00000000000000000000000000000010;
REG[59] <= 32'b00000000000000000000000000000000;
REG[60] <= 32'b00000000000000000000000000000000;
REG[61] <= 32'b00000000000000000000000000000000;
REG[62] <= 32'b00000000000000000000000000000000;
REG[63] <= 32'b00000000000000000000000000000000;
REG[64] <= 32'b00000000000101000000001100000000;
REG[65] <= 32'b00000000000000000000000000000000;
REG[66] <= 32'b00000000000001000000000000000000;
REG[67] <= 32'b00000000000000000000000000000000;
REG[68] <= 32'b00000000000000000000000000001111;
REG[69] <= 32'b00000101000110100000110100000000;
REG[70] <= 32'b00000000000000000000000000000000;
REG[71] <= 32'b00001011000000000000000000000000;
REG[72] <= 32'b00000000000000000000000000000000;
REG[73] <= 32'b00000000000000000000000000000000;
REG[74] <= 32'b00000000000000000000000000000000;
REG[75] <= 32'b00000000000011000001010000000000;
REG[76] <= 32'b00001000000000000000000000011011;
REG[77] <= 32'b00001001000000000000000000000000;
REG[78] <= 32'b00000000000000000000000000000000;
REG[79] <= 32'b00101001001111110000000000000000;
REG[80] <= 32'b00000000000000000000000000000000;
REG[81] <= 32'b00000000000000000000000000000000;
REG[82] <= 32'b00000011001010010000000000000000;
REG[83] <= 32'b00000000000000000000000100000000;
REG[84] <= 32'b00000000000000000000000000000000;
REG[85] <= 32'b00000000000000000000000000000000;
REG[86] <= 32'b00000000000000000000000000000000;
REG[87] <= 32'b00000101000000000000000000000000;
REG[88] <= 32'b00000000000000110000000000000000;
REG[89] <= 32'b00000000000000000000000000000000;
REG[90] <= 32'b00000000000000000000000000001001;
REG[91] <= 32'b00000000000000000000001000001100;
REG[92] <= 32'b00000000000000000000000000000000;
REG[93] <= 32'b00000000000000000000000000100010;
REG[94] <= 32'b00000000000000000000001100010110;
REG[95] <= 32'b00010001000000000000000000000000;
REG[96] <= 32'b00000000000000000000000000000000;
REG[97] <= 32'b00000000000000000000000000000000;
REG[98] <= 32'b00000000000000000000000000000000;
REG[99] <= 32'b00000000000000000000000000000000;
REG[100] <= 32'b00010011000000000000000000010100;
REG[101] <= 32'b00000011000000000000000000000000;
REG[102] <= 32'b00000000000000000000000000000000;
REG[103] <= 32'b00000000000000000000000000011000;
REG[104] <= 32'b00000000000000000000000000000000;
REG[105] <= 32'b00000000000000000000000000000000;
REG[106] <= 32'b00000000000000000000000000000000;
REG[107] <= 32'b00000000000000000000000000000000;
REG[108] <= 32'b00000000000000000000000000000000;
REG[109] <= 32'b00000000000000000000000000000000;
REG[110] <= 32'b00000000000000000000000000000000;
REG[111] <= 32'b00000000000000000000000000000000;
REG[112] <= 32'b00000100000000000000000000000000;
REG[113] <= 32'b00000000000000000000000000011011;
REG[114] <= 32'b00000000000000000000000000000000;
REG[115] <= 32'b00010100000000000000000000000000;
REG[116] <= 32'b00000000000000000000000000000100;
REG[117] <= 32'b00000000000000000000000000000000;
REG[118] <= 32'b00000000000000000000000000000000;
REG[119] <= 32'b00000000000000000000000000000000;
REG[120] <= 32'b00000000000000000000000000000000;
REG[121] <= 32'b00000000000000000000000000000000;
REG[122] <= 32'b00000000000000000000000000000000;
REG[123] <= 32'b00000000000110010000000000000000;
REG[124] <= 32'b00000000000000000000000000011100;
REG[125] <= 32'b00000000000000000000000000000000;
REG[126] <= 32'b00000000000101100000000000000000;
REG[127] <= 32'b00000000000000000000000000000000;
REG[128] <= 32'b00000000000000000000000000000000;
REG[129] <= 32'b00000000000011100000000000000000;
REG[130] <= 32'b00000000000000000000000000000000;
REG[131] <= 32'b00000000000000000000000000000000;
REG[132] <= 32'b00000000000000000000000000000000;
REG[133] <= 32'b00000000000000000000000000000000;
REG[134] <= 32'b00000000000000000000000000000000;
REG[135] <= 32'b00001001001101010001110100000000;
REG[136] <= 32'b00000000000000000000000000000111;
REG[137] <= 32'b01000100000000000000000000000000;
REG[138] <= 32'b00000000000101110000011100000000;
REG[139] <= 32'b00000000000000000000000000000000;
REG[140] <= 32'b00000111000000000000000000000000;
REG[141] <= 32'b00000000000000000000010000000000;
REG[142] <= 32'b00000000000000000000000000000000;
REG[143] <= 32'b00000000000000000000000000000000;
REG[144] <= 32'b00000000000000000000000000000000;
REG[145] <= 32'b00000000000000000000000000000000;
REG[146] <= 32'b00000000000000000000000000000000;
REG[147] <= 32'b00000000000000110010001000000000;
REG[148] <= 32'b00000000000000100000000000000000;
REG[149] <= 32'b00000000000000000111111100101111;
REG[150] <= 32'b00000000000000000000000000000000;
REG[151] <= 32'b00000000000000000000000000010101;
REG[152] <= 32'b00000000000000000101010100000000;
REG[153] <= 32'b00000000000000000000000000000000;
REG[154] <= 32'b00001111000000000000000000011101;
REG[155] <= 32'b00000000000000000100011000000000;
REG[156] <= 32'b00000000000000000000000000000000;
REG[157] <= 32'b00000000000000000000000000000000;
REG[158] <= 32'b00000000000000000000000000000000;
REG[159] <= 32'b00101010000001110000000000000000;
REG[160] <= 32'b00000001000011000001110100101110;
REG[161] <= 32'b00000000001010110100000101011011;
REG[162] <= 32'b00000000000000000000000000000000;
REG[163] <= 32'b00001001000000100000000000001111;
REG[164] <= 32'b00000111000000000000000000000000;
REG[165] <= 32'b00000000000000000000000000000000;
REG[166] <= 32'b00000000000001000000000000000000;
REG[167] <= 32'b00001101000000000000000000000000;
REG[168] <= 32'b00000000000000000000000000000000;
REG[169] <= 32'b00000000000000000000000000000000;
REG[170] <= 32'b00000000000000000000000000000000;
REG[171] <= 32'b00000000000011110000000000000000;
REG[172] <= 32'b00000000000000000000000000010011;
REG[173] <= 32'b00000000000000000000001100001011;
REG[174] <= 32'b00000000000000000000000000000000;
REG[175] <= 32'b00000000000000000000000000111010;
REG[176] <= 32'b00000000000000000000000100000110;
REG[177] <= 32'b00000000000000010000000000000000;
REG[178] <= 32'b00000000000000000000000000101010;
REG[179] <= 32'b00000000000000000001110100000000;
REG[180] <= 32'b00000000000000000000000000000000;
REG[181] <= 32'b00000000000000000000000000000000;
REG[182] <= 32'b00000000000000000000000000000000;
REG[183] <= 32'b00011011001110010000110000000000;
REG[184] <= 32'b00000000000000000000000000000000;
REG[185] <= 32'b00000000001101010001100100000000;
REG[186] <= 32'b00000000000000000000000000000000;
REG[187] <= 32'b00000000000000000000000000000000;
REG[188] <= 32'b00000000000100010000000000000100;
REG[189] <= 32'b00000000000000000000000000000000;
REG[190] <= 32'b00000000000000000000000000000000;
REG[191] <= 32'b00000000000000000000000000010010;
REG[192] <= 32'b00000000000000000000000000000000;
REG[193] <= 32'b00000000000000000000000000000000;
REG[194] <= 32'b00000000000000000000000000000000;
REG[195] <= 32'b00000000000000000000000000000000;
REG[196] <= 32'b00001101000111000000000000000000;
REG[197] <= 32'b00000000000000000011010000000110;
REG[198] <= 32'b00000000000000000000000000000000;
REG[199] <= 32'b00010100000000000000000000000000;
REG[200] <= 32'b00000000000000000010101100000000;
REG[201] <= 32'b00000000000001100000000000000000;
REG[202] <= 32'b00101101000010110000000000000000;
REG[203] <= 32'b00000000000000000010010100000000;
REG[204] <= 32'b00000000000000000000000000000000;
REG[205] <= 32'b00000000000000000000000000000000;
REG[206] <= 32'b00000000000000000000000000000000;
REG[207] <= 32'b00000000000000000000000000001101;
REG[208] <= 32'b00010000000110000000000000000000;
REG[209] <= 32'b00000000000000000001010100110011;
REG[210] <= 32'b00000000000000000000000000000000;
REG[211] <= 32'b00010101000011100000000000000000;
REG[212] <= 32'b00000000000000000000000000011011;
REG[213] <= 32'b00000000000000000000000000000000;
REG[214] <= 32'b00001010000011000000000000000000;
REG[215] <= 32'b00000000000000000000000000000000;
REG[216] <= 32'b00000000000000000000000000000000;
REG[217] <= 32'b00000000000000000000000000000000;
REG[218] <= 32'b00000000000000000000000000000000;
REG[219] <= 32'b00000000000000000000000000000000;
REG[220] <= 32'b00010100000000000000000000000000;
REG[221] <= 32'b00000000000000000011001000000000;
REG[222] <= 32'b00000000001011000000000000000000;
REG[223] <= 32'b00000100000000000000000000000000;
REG[224] <= 32'b00000000000000000000100000000000;
REG[225] <= 32'b00000000010010000000000000000000;
REG[226] <= 32'b00000000000000000000000000000000;
REG[227] <= 32'b00001001000000000000000000000000;
REG[228] <= 32'b00000000000000000000000000000000;
REG[229] <= 32'b00000000000000000000000000000000;
REG[230] <= 32'b00000000000000000000000000000000;
REG[231] <= 32'b00000000000000000000000000000000;
REG[232] <= 32'b00000000000011000000000000000000;
REG[233] <= 32'b00000000000000000000000000000011;
REG[234] <= 32'b00011000001011100010100100000000;
REG[235] <= 32'b00000001000010110000000000000000;
REG[236] <= 32'b00000000000000000000100000000000;
REG[237] <= 32'b00000000000100010010000000000000;
REG[238] <= 32'b00000000000011010000000000000000;
REG[239] <= 32'b00000000000000000000000000010100;
REG[240] <= 32'b00000000000000000000000000000000;
REG[241] <= 32'b00000000000000000000000000000000;
REG[242] <= 32'b00000000000000000000000000000000;
REG[243] <= 32'b00000000000000000000000000000000;
REG[244] <= 32'b00000000000000000000000000000000;
REG[245] <= 32'b00000000000000000000000000000000;
REG[246] <= 32'b00000000000000000000000000000000;
REG[247] <= 32'b00000000000000000000000000000000;
REG[248] <= 32'b00001101000000000000011100000000;
REG[249] <= 32'b00000000001100010001111100000000;
REG[250] <= 32'b00000000000000000000000000000000;
REG[251] <= 32'b00100010000000000000000000000000;
REG[252] <= 32'b00000000000000000000000000000000;
REG[253] <= 32'b00000000000000000000000000000000;
REG[254] <= 32'b00000000000000000000000000000000;
REG[255] <= 32'b00000000000000000000000000000000;
REG[256] <= 32'b00010101000000110000000000000000;
REG[257] <= 32'b00000000000000000000000000000000;
REG[258] <= 32'b00000000000000000000000000000000;
REG[259] <= 32'b00001011000000000000110100000000;
REG[260] <= 32'b00000000000000000000000000000000;
REG[261] <= 32'b00000000000000000000000000000000;
REG[262] <= 32'b00000000000000000100010000000000;
REG[263] <= 32'b00000000000000000000000000000000;
REG[264] <= 32'b00000000000000000000000000000000;
REG[265] <= 32'b00000000000000000000000000000000;
REG[266] <= 32'b00000000000000000000000000000000;
REG[267] <= 32'b00000000000010000000000000000000;
REG[268] <= 32'b00000000000000010000000000000010;
REG[269] <= 32'b00000000000000000000111100010011;
REG[270] <= 32'b00000000000101110000000000000000;
REG[271] <= 32'b00000000000000000000000000010111;
REG[272] <= 32'b00001111000000000000010100000000;
REG[273] <= 32'b00000000000100000000000000000000;
REG[274] <= 32'b00000000000000000000000000100110;
REG[275] <= 32'b00001110000000000000000000000000;
REG[276] <= 32'b00000000000000000000000000000000;
REG[277] <= 32'b00000000000000000000000000000000;
REG[278] <= 32'b00000000000000000000000000000000;
REG[279] <= 32'b00000000000000000000000000001000;
REG[280] <= 32'b00000000000000000000000000000000;
REG[281] <= 32'b00000000000101000001011000010111;
REG[282] <= 32'b00000000000000000000000000001110;
REG[283] <= 32'b00000000000000000000000000000000;
REG[284] <= 32'b00000000000010100001110100011101;
REG[285] <= 32'b00000000000000000000000000010001;
REG[286] <= 32'b00000000000000000000000000000000;
REG[287] <= 32'b00000000000010010010001000011011;
REG[288] <= 32'b00000000000000000000000000000000;
REG[289] <= 32'b00000000000000000000000000000000;
REG[290] <= 32'b00000000000000000000000000000000;
REG[291] <= 32'b00000000000000000000000000000000;
REG[292] <= 32'b00000000000000000000000000000000;
REG[293] <= 32'b00000000000000000001010100000010;
REG[294] <= 32'b00000000000000000000000000000000;
REG[295] <= 32'b00000000000000000000000000000000;
REG[296] <= 32'b00000000000000000000000000000000;
REG[297] <= 32'b00000000000000000000000000000000;
REG[298] <= 32'b00000000000000000000000000000000;
REG[299] <= 32'b00000000000000000000010100000000;
REG[300] <= 32'b00000000000000000000000000000000;
REG[301] <= 32'b00000000000000000000000000000000;
REG[302] <= 32'b00000000000000000000000000000000;
REG[303] <= 32'b00000000000000000000000000001100;
REG[304] <= 32'b00010010000011010000000000010010;
REG[305] <= 32'b00000000001000110011000100010111;
REG[306] <= 32'b00000000000001000000000000000000;
REG[307] <= 32'b00001000000001100000000000000000;
REG[308] <= 32'b00000000000001010011000100000100;
REG[309] <= 32'b00000000000000000000001000000000;
REG[310] <= 32'b00011000000011010000000000000000;
REG[311] <= 32'b00000000000000000000000000010010;
REG[312] <= 32'b00000000000000000000000000000000;
REG[313] <= 32'b00000000000000000000000000000000;
REG[314] <= 32'b00000000000000000000000000000000;
REG[315] <= 32'b00000000000110010000000000000000;
REG[316] <= 32'b00000000000000000000000000000110;
REG[317] <= 32'b00000000000000000000000000000000;
REG[318] <= 32'b00000000001010100000110000000000;
REG[319] <= 32'b00000000000000000000000000010010;
REG[320] <= 32'b00000000000000000000000000000000;
REG[321] <= 32'b00000000000111010000011100000000;
REG[322] <= 32'b00000000000000000000000000001000;
REG[323] <= 32'b00000000000000000000000000000000;
REG[324] <= 32'b00000000000000000000000000000000;
REG[325] <= 32'b00000000000000000000000000000000;
REG[326] <= 32'b00000000000000000000000000000000;
REG[327] <= 32'b00000000000000000000000000000000;
REG[328] <= 32'b00000000000000000000011100001001;
REG[329] <= 32'b00000000000000000000000000000000;
REG[330] <= 32'b00000000000000000000000000000000;
REG[331] <= 32'b00000000000000000000000000001111;
REG[332] <= 32'b00000101000001000000111000000000;
REG[333] <= 32'b00000000000000000000000000000000;
REG[334] <= 32'b00000000000000000000000000000000;
REG[335] <= 32'b00000000000000000000100000000000;
REG[336] <= 32'b00000000000000000000000000000000;
REG[337] <= 32'b00000000000000000000000000000000;
REG[338] <= 32'b00000000000000000000000000000000;
REG[339] <= 32'b00000000000000000001000000000000;
REG[340] <= 32'b00000000000000000000000000100111;
REG[341] <= 32'b00010010000000000000000000000000;
REG[342] <= 32'b00000000000000000001011000000000;
REG[343] <= 32'b00000011000000000000000000011101;
REG[344] <= 32'b00000000000000000000000000001000;
REG[345] <= 32'b00000000000000000000111000000000;
REG[346] <= 32'b00100010000000000000000000000000;
REG[347] <= 32'b00000000000000000000000000010001;
REG[348] <= 32'b00000000000000000000000000000000;
REG[349] <= 32'b00000000000000000000000000000000;
REG[350] <= 32'b00000000000000000000000000000000;
REG[351] <= 32'b00000000000000000000000000000000;
REG[352] <= 32'b00000000000000000000000000000000;
REG[353] <= 32'b00000000000000000010000000010101;
REG[354] <= 32'b00010001000000000000000000000000;
REG[355] <= 32'b00000000000000000000000000000000;
REG[356] <= 32'b00000000000000000000000000000000;
REG[357] <= 32'b00011110000000000000000000000000;
REG[358] <= 32'b00000000000000000000000000000000;
REG[359] <= 32'b00000000000001000000000000000001;
REG[360] <= 32'b00000000000000000000000000000000;
REG[361] <= 32'b00000000000000000000000000000000;
REG[362] <= 32'b00000000000000000000000000000000;
REG[363] <= 32'b00000000000000000000000000000000;
REG[364] <= 32'b00101010001001100000000000001000;
REG[365] <= 32'b01010101000000000000000000000000;
REG[366] <= 32'b00000000000010010000000000000000;
REG[367] <= 32'b00101000000010110000000000000000;
REG[368] <= 32'b00010001000000000000000000000000;
REG[369] <= 32'b00000000000110000000000000000000;
REG[370] <= 32'b00011100000000110000000000000000;
REG[371] <= 32'b01000000000000000000000000001010;
REG[372] <= 32'b00000000000000000000000000000000;
REG[373] <= 32'b00000000000000000000000000000000;
REG[374] <= 32'b00000000000000000000000000000000;
REG[375] <= 32'b00000000000000000000000000000000;
REG[376] <= 32'b00000000000000000110000100011111;
REG[377] <= 32'b00110100000110010001011000000000;
REG[378] <= 32'b00000000000011110001000100000000;
REG[379] <= 32'b00000000000000000010010100000000;
REG[380] <= 32'b00000000000000000000000000000000;
REG[381] <= 32'b00000000000000000000001100000000;
REG[382] <= 32'b00000000000000000010111100000000;
REG[383] <= 32'b00000000000001110000000000000000;
REG[384] <= 32'b00000000000000000000000000000000;
REG[385] <= 32'b00000000000000000000000000000000;
REG[386] <= 32'b00000000000000000000000000000000;
REG[387] <= 32'b00000000001011000000000000000000;
REG[388] <= 32'b00000000000000000000000000000000;
REG[389] <= 32'b00000000000000000010111000110111;
REG[390] <= 32'b00000000001100100000000000000000;
REG[391] <= 32'b00000000000000000000000000000000;
REG[392] <= 32'b00000000000000000001100100000000;
REG[393] <= 32'b00000000001100010000000000000000;
REG[394] <= 32'b00000000000000000000000000100010;
REG[395] <= 32'b00100000000000000010010100010011;
REG[396] <= 32'b00000000000000000000000000000000;
REG[397] <= 32'b00000000000000000000000000000000;
REG[398] <= 32'b00000000000000000000000000000000;
REG[399] <= 32'b00000000000100010001000000000000;
REG[400] <= 32'b00000000000000000000000000000000;
REG[401] <= 32'b00000000001111100001001100000101;
REG[402] <= 32'b00000000000000000000000000000000;
REG[403] <= 32'b00000000000000000000000000000000;
REG[404] <= 32'b00000000000000110000101000000000;
REG[405] <= 32'b00000000000000000000000000000000;
REG[406] <= 32'b00000000000000000000000100000000;
REG[407] <= 32'b00000000000011000000100100000000;
REG[408] <= 32'b00000000000000000000000000000000;
REG[409] <= 32'b00000000000000000000000000000000;
REG[410] <= 32'b00000000000000000000000000000000;
REG[411] <= 32'b00000000000000000000000000000000;
REG[412] <= 32'b00000000000110000000000000000000;
REG[413] <= 32'b00000000000000000010011000100110;
REG[414] <= 32'b00000000000000000000000000000000;
REG[415] <= 32'b00000000000000000000000000000000;
REG[416] <= 32'b00000000000000000010011100010000;
REG[417] <= 32'b00000000000000000000000000000000;
REG[418] <= 32'b00000000000000000000000000110110;
REG[419] <= 32'b00100101000000000000110100000000;
REG[420] <= 32'b00000000000000000000000000000000;
REG[421] <= 32'b00000000000000000000000000000000;
REG[422] <= 32'b00000000000000000000000000000000;
REG[423] <= 32'b00000000000000000000000000001001;
REG[424] <= 32'b00000000000000000011011100101000;
REG[425] <= 32'b00000000000011100000000000000000;
REG[426] <= 32'b00000001000101010000000000000000;
REG[427] <= 32'b00000000000000000010010000000110;
REG[428] <= 32'b00000000000011010000100100000000;
REG[429] <= 32'b00000000000100000000000000000000;
REG[430] <= 32'b00000000000000000010010000010010;
REG[431] <= 32'b00000110000000000001111100000000;
REG[432] <= 32'b00000000000000000000000000000000;
REG[433] <= 32'b00000000000000000000000000000000;
REG[434] <= 32'b00000000000000000000000000000000;
REG[435] <= 32'b00000000000000000000010100000000;
REG[436] <= 32'b00000000000000000000000000000000;
REG[437] <= 32'b00000101000000000000000000000000;
REG[438] <= 32'b00000000000000000000000000000000;
REG[439] <= 32'b00000000000000000000000000000000;
REG[440] <= 32'b00000000000000000000100100010011;
REG[441] <= 32'b00000000000000000000000000000000;
REG[442] <= 32'b00000000000000000000000000000000;
REG[443] <= 32'b00000000000000000000000000000000;
REG[444] <= 32'b00000000000000000000000000000000;
REG[445] <= 32'b00000000000000000000000000000000;
REG[446] <= 32'b00000000000000000000000000000000;
REG[447] <= 32'b00000000000000000000000000000000;
REG[448] <= 32'b00000000000000000000000000000000;
REG[449] <= 32'b00000000000000000000000000000000;
REG[450] <= 32'b00000000000000000000000000000000;
REG[451] <= 32'b00000110000000000000000000000000;
REG[452] <= 32'b00000000000010110000000000000000;
REG[453] <= 32'b00000000000000000000000000000000;
REG[454] <= 32'b00001111000000000000000000000000;
REG[455] <= 32'b00000000000000100000000000000000;
REG[456] <= 32'b00000000000000000000000000000000;
REG[457] <= 32'b00000000000000000000000000000000;
REG[458] <= 32'b00000000000000000000000000000000;
REG[459] <= 32'b00000000000000000000000000000000;
REG[460] <= 32'b00000000000000000000000000000000;
REG[461] <= 32'b00000000000000000001101100000000;
REG[462] <= 32'b00000000000000000000000000000000;
REG[463] <= 32'b00000000000000000000000000000000;
REG[464] <= 32'b00000111000000000000000000000000;
REG[465] <= 32'b00000000000001000000000000000000;
REG[466] <= 32'b00000000000000000000000000000000;
REG[467] <= 32'b00010000000000000001100100000000;
REG[468] <= 32'b00000000000000000000000000000000;
REG[469] <= 32'b00000000000000000000000000000000;
REG[470] <= 32'b00000000000000000000000000000000;
REG[471] <= 32'b00000000000000000000000000000000;
REG[472] <= 32'b00000000000000000000000000011110;
REG[473] <= 32'b00010010000000000000011100001101;
REG[474] <= 32'b00000000000000000000000000000000;
REG[475] <= 32'b00000000000000000000000000000000;
REG[476] <= 32'b00000000000000000000000000000000;
REG[477] <= 32'b00000000000000000000000000000000;
REG[478] <= 32'b00000000000000000000000000000000;
REG[479] <= 32'b00000000000000000000000000010011;
REG[480] <= 32'b00000000000000000000000000000000;
REG[481] <= 32'b00000000000000000000000000000000;
REG[482] <= 32'b00000000000000000000000000000000;
REG[483] <= 32'b00000000000000000000010000000000;
REG[484] <= 32'b00000000000000000000000000000000;
REG[485] <= 32'b00000011000000000000000000000000;
REG[486] <= 32'b00000000000000000000000000000000;
REG[487] <= 32'b00000000000000000000000000000000;
REG[488] <= 32'b00000000000000000000000000000000;
REG[489] <= 32'b00000000000000000000000000000000;
REG[490] <= 32'b00000000000110110000000000000000;
REG[491] <= 32'b00010101000000000000000000000000;
REG[492] <= 32'b00000000000000000000000000000000;
REG[493] <= 32'b00000000000000000000000000000000;
REG[494] <= 32'b00000000000000000000000000000000;
REG[495] <= 32'b00000000000000000000000000011000;
REG[496] <= 32'b00010010000000000010000100101011;
REG[497] <= 32'b00011101000000000001111000000000;
REG[498] <= 32'b00000000000000000000000000010010;
REG[499] <= 32'b00000000000000000000000000000000;
REG[500] <= 32'b00100010000000000001100100000000;
REG[501] <= 32'b00000000000000000000000000100000;
REG[502] <= 32'b00000000000000000000111100001000;
REG[503] <= 32'b00010001000000000001110000000010;
REG[504] <= 32'b00000000000000000000000000000000;
REG[505] <= 32'b00000000000000000000000000000000;
REG[506] <= 32'b00000000000000000000000000000000;
REG[507] <= 32'b00000000000001010000100000000000;
REG[508] <= 32'b00000000000000000000000000000000;
REG[509] <= 32'b00000000000000000000000000000000;
REG[510] <= 32'b00000000000000000000111100000000;
REG[511] <= 32'b00000000000000000000000000001011;
REG[512] <= 32'b00000000000000000000000000000000;
REG[513] <= 32'b00000000000000000000000000000000;
REG[514] <= 32'b00000000000000000000000000010010;
REG[515] <= 32'b00000000000000000000000000001011;
REG[516] <= 32'b00000000000000000000000000000000;
REG[517] <= 32'b00000000000000000000000000000000;
REG[518] <= 32'b00000000000000000000000000000000;
REG[519] <= 32'b00000100000000000000010000000000;
REG[520] <= 32'b00000000000000000000000000000000;
REG[521] <= 32'b00000000000010010000000100000000;
REG[522] <= 32'b00011111001100110100001100000000;
REG[523] <= 32'b00000000000000000000000000000000;
REG[524] <= 32'b00000000000000000000000000000000;
REG[525] <= 32'b00010010001101100011011000000000;
REG[526] <= 32'b00000000000000000000000000000000;
REG[527] <= 32'b00000000000010000000000000000000;
REG[528] <= 32'b00000000000000000000000000000000;
REG[529] <= 32'b00000000000000000000000000000000;
REG[530] <= 32'b00000000000000000000000000000000;
REG[531] <= 32'b00000000000000000000000000000000;
REG[532] <= 32'b00001100000000000000000000000000;
REG[533] <= 32'b00000000000000000000001000110110;
REG[534] <= 32'b00000000000000000000000000000000;
REG[535] <= 32'b00100000000111100000000000000000;
REG[536] <= 32'b00000000000000000000000000000000;
REG[537] <= 32'b00000000000000000000000000000000;
REG[538] <= 32'b00000000001000110000000000000100;
REG[539] <= 32'b00000000000000000000000000000000;
REG[540] <= 32'b00000000000000000000000000000000;
REG[541] <= 32'b00000000000000000000000000000000;
REG[542] <= 32'b00000000000000000000000000000000;
REG[543] <= 32'b00000000000000000000000000001100;
REG[544] <= 32'b00011110001110000000000000000110;
REG[545] <= 32'b00000000001000000000000000000000;
REG[546] <= 32'b00000000000000000000000000100010;
REG[547] <= 32'b00000000000111000000000000000000;
REG[548] <= 32'b00000000000000000000011100000000;
REG[549] <= 32'b00000000000000000000000001010110;
REG[550] <= 32'b00000110000000000000000000000000;
REG[551] <= 32'b00000000000000000000000000000000;
REG[552] <= 32'b00000000000000000000000000000000;
REG[553] <= 32'b00000000000000000000000000000000;
REG[554] <= 32'b00000000000000000000000000000000;
REG[555] <= 32'b00000000000000000000000000000000;
REG[556] <= 32'b00000000000000000000000000011101;
REG[557] <= 32'b00000000000000000000000000000000;
REG[558] <= 32'b00000000000000000000000000000000;
REG[559] <= 32'b00000000000000000000000000011111;
REG[560] <= 32'b00010101000000000000000000000000;
REG[561] <= 32'b00000000000000000000000000000000;
REG[562] <= 32'b00000000000000000000000000000000;
REG[563] <= 32'b00000000000000000000000000000000;
REG[564] <= 32'b00000000000000000000000000000000;
REG[565] <= 32'b00000000000000000000000000000000;
REG[566] <= 32'b00000000000000000000000000000000;
REG[567] <= 32'b00001110000000000000000000010010;
REG[568] <= 32'b00010110000100110000000000000000;
REG[569] <= 32'b00000101000000000000000000000000;
REG[570] <= 32'b00000010000000000000000000000000;
REG[571] <= 32'b00000111000010110000000000000000;
REG[572] <= 32'b00001110000000000000000000001011;
REG[573] <= 32'b00001011000000000000000000000000;
REG[574] <= 32'b00000000000000000000000000000000;
REG[575] <= 32'b00000000000000000000001100010010;
REG[576] <= 32'b00000000000000000000000000000000;
REG[577] <= 32'b00000000000000000000000000000000;
REG[578] <= 32'b00000000000000000000000000000000;
REG[579] <= 32'b00000000000000100000001100000000;
REG[580] <= 32'b00000011000000000000000000000000;
REG[581] <= 32'b00000000000000000001100100010001;
REG[582] <= 32'b00000000000000000000000000000000;
REG[583] <= 32'b00010010000000000000000000000000;
REG[584] <= 32'b00000000000000000000000000000000;
REG[585] <= 32'b00000000000000000000000000000000;
REG[586] <= 32'b00011110000000000000000000000000;
REG[587] <= 32'b00000000000000000000110000000000;
REG[588] <= 32'b00000000000000000000000000000000;
REG[589] <= 32'b00000000000000000000000000000000;
REG[590] <= 32'b00000000000000000000000000000000;
REG[591] <= 32'b00000000000000000000000000000000;
REG[592] <= 32'b00000000000000000001100100001110;
REG[593] <= 32'b00000000000010000000000000010010;
REG[594] <= 32'b00001001000000000000000000000000;
REG[595] <= 32'b00000000000000000000100000001100;
REG[596] <= 32'b00000000000000000000000000010100;
REG[597] <= 32'b00001101000101000000011100000000;
REG[598] <= 32'b00000000000000000000000000011110;
REG[599] <= 32'b00110000000000000000000100001100;
REG[600] <= 32'b00000000000000000000000000000000;
REG[601] <= 32'b00000000000000000000000000000000;
REG[602] <= 32'b00000000000000000000000000000000;
REG[603] <= 32'b00000000000000000001111000000000;
REG[604] <= 32'b00000010000001010000000000000000;
REG[605] <= 32'b00000000000000000001110000000000;
REG[606] <= 32'b00000000000000000000001000000000;
REG[607] <= 32'b00000000000000000000000000011000;
REG[608] <= 32'b00100000000000000000111000000000;
REG[609] <= 32'b00000000000000000000000000000000;
REG[610] <= 32'b00000000000000000000000000001111;
REG[611] <= 32'b00001100000000000000000000000000;
REG[612] <= 32'b00000000000000000000000000000000;
REG[613] <= 32'b00000000000000000000000000000000;
REG[614] <= 32'b00000000000000000000000000000000;
REG[615] <= 32'b00101101000000000000000000000000;
REG[616] <= 32'b00000000000000000000000000000000;
REG[617] <= 32'b00000000000000000011100100111101;
REG[618] <= 32'b00100010000000000000000000000000;
REG[619] <= 32'b00000111000000000000011100000000;
REG[620] <= 32'b00000000000000000000011000001110;
REG[621] <= 32'b00000000000000000000000000000000;
REG[622] <= 32'b00000000000000000000000000000000;
REG[623] <= 32'b00000000000000000000000000000000;
REG[624] <= 32'b00000000000000000000000000000000;
REG[625] <= 32'b00000000000000000000000000000000;
REG[626] <= 32'b00000000000000000000000000000000;
REG[627] <= 32'b00000000001010110000000000000000;
REG[628] <= 32'b00000000000000000000000000000000;
REG[629] <= 32'b00000000000000000000100000000000;
REG[630] <= 32'b00000000001110110000011100000000;
REG[631] <= 32'b00000000000000000000000000011001;
REG[632] <= 32'b00000000000000000000001000000000;
REG[633] <= 32'b00000000000100000010101100000000;
REG[634] <= 32'b00000000000000000000000000000000;
REG[635] <= 32'b00000000000000000000000000000000;
REG[636] <= 32'b00000000000000000000000000000000;
REG[637] <= 32'b00000000000000000000000000000000;
REG[638] <= 32'b00000000000000000000000000000000;
REG[639] <= 32'b00000000000110010011101100000000;
REG[640] <= 32'b00000000000000000001000000101100;
REG[641] <= 32'b00000000000001000000101000000110;
REG[642] <= 32'b00000000000000000010000000000000;
REG[643] <= 32'b00000000000000000000000000011100;
REG[644] <= 32'b00011000000000000000000100010100;
REG[645] <= 32'b00001101000000000000000000000000;
REG[646] <= 32'b00000000000000000000000000000000;
REG[647] <= 32'b00001000000000000000000000010011;
REG[648] <= 32'b00000000000000000000000000000000;
REG[649] <= 32'b00000000000000000000000000000000;
REG[650] <= 32'b00000000000000000000000000000000;
REG[651] <= 32'b00000000000000000000000000000000;
REG[652] <= 32'b00000000000000000000000000000000;
REG[653] <= 32'b00001000000000000001100000011011;
REG[654] <= 32'b00000000000000000000000000000000;
REG[655] <= 32'b00010100000000000000000000000000;
REG[656] <= 32'b00000000000000000001100100000000;
REG[657] <= 32'b00000000000101000000000000000000;
REG[658] <= 32'b00000000000001000000000000000000;
REG[659] <= 32'b00000000000000000010101000000000;
REG[660] <= 32'b00000000000000000000000000000000;
REG[661] <= 32'b00000000000000000000000000000000;
REG[662] <= 32'b00000000000000000000000000000000;
REG[663] <= 32'b00000000000000000000000000000000;
REG[664] <= 32'b00001011001011010000000000000000;
REG[665] <= 32'b00000000000100000000000000000000;
REG[666] <= 32'b00000000000000000000000000000000;
REG[667] <= 32'b00000000000111000000000000000000;
REG[668] <= 32'b00000000000000000000000000000000;
REG[669] <= 32'b00000000000000000000000000000000;
REG[670] <= 32'b00000000000000000000000000000000;
REG[671] <= 32'b00000000000000000000000000000000;
REG[672] <= 32'b00000000000000000000000000000000;
REG[673] <= 32'b00000000000000000000000000000000;
REG[674] <= 32'b00000000000000000000000000000000;
REG[675] <= 32'b00000000000000000001110000000000;
REG[676] <= 32'b00000000000000000000000000000000;
REG[677] <= 32'b00000000000000000000000000001010;
REG[678] <= 32'b00000000000000000000000000000000;
REG[679] <= 32'b00001000000000000000000000000000;
REG[680] <= 32'b00000000000000000000000000000000;
REG[681] <= 32'b00000000000000000000000000000000;
REG[682] <= 32'b00000000000000000000000000000000;
REG[683] <= 32'b00000000000000000000000000000000;
REG[684] <= 32'b00000000000000000000000000000000;
REG[685] <= 32'b00000000000000000000000000000000;
REG[686] <= 32'b00000000000000000000000000000000;
REG[687] <= 32'b00100000000000000000000000000000;
REG[688] <= 32'b00000000000000000000000000000000;
REG[689] <= 32'b00000000000011000000000000000000;
REG[690] <= 32'b00101001000000000000000000000000;
REG[691] <= 32'b00000000000000000000000000000000;
REG[692] <= 32'b00000000000000000000000000000000;
REG[693] <= 32'b00110001001100110000000000000000;
REG[694] <= 32'b00000000000000000000000000000000;
REG[695] <= 32'b00000000000000000000000000000000;
REG[696] <= 32'b00000000000000000000000000000000;
REG[697] <= 32'b00000000000000000000000000000000;
REG[698] <= 32'b00000000000000000000000000000000;
REG[699] <= 32'b00000000001111010011010100000000;
REG[700] <= 32'b00001011000010000000000000000000;
REG[701] <= 32'b00000000000000000010110100001001;
REG[702] <= 32'b00000000000001000000000000000000;
REG[703] <= 32'b00000000000000000000000000000000;
REG[704] <= 32'b00000000000000000000000000000000;
REG[705] <= 32'b00000000000101000000001100000000;
REG[706] <= 32'b00000000000000000000000000000000;
REG[707] <= 32'b00000000000000000000000000000111;
REG[708] <= 32'b00000000000000000000000000000000;
REG[709] <= 32'b00000000000000000000000000000000;
REG[710] <= 32'b00000000000000000000000000000000;
REG[711] <= 32'b00010100000011010010101000000100;
REG[712] <= 32'b00001000000000000000000000000000;
REG[713] <= 32'b00000000000000000000100001000100;
REG[714] <= 32'b00000000000000000000000100000000;
REG[715] <= 32'b00001011000000000011100101111111;
REG[716] <= 32'b01000011000000000000000000000000;
REG[717] <= 32'b00000000000000000000000000000000;
REG[718] <= 32'b00011000000100110000000001000111;
REG[719] <= 32'b01000100000010110000000000000000;
REG[720] <= 32'b00000000000000000000000000000000;
REG[721] <= 32'b00000000000000000000000000000000;
REG[722] <= 32'b00000000000000000000000000000000;
REG[723] <= 32'b00000000000000000000000000000000;
REG[724] <= 32'b00100100001000110000000000000001;
REG[725] <= 32'b00011011000000000000000000000000;
REG[726] <= 32'b00000000000000000000000000000000;
REG[727] <= 32'b00110111000000000000000000000000;
REG[728] <= 32'b00000000000000000000000000000000;
REG[729] <= 32'b00000000000000000000000000000000;
REG[730] <= 32'b00010011000000000000000000000000;
REG[731] <= 32'b00000000000000000001000100000000;
REG[732] <= 32'b00000000000000000000000000000000;
REG[733] <= 32'b00000000000000000000000000000000;
REG[734] <= 32'b00000000000000000000000000000000;
REG[735] <= 32'b00000000000000000000000000001100;
REG[736] <= 32'b00001000000000000000000000000000;
REG[737] <= 32'b00000000000000000000000000000000;
REG[738] <= 32'b00000000000000000000000000000000;
REG[739] <= 32'b00000000000000000000000000011000;
REG[740] <= 32'b00001100000000000000000000000000;
REG[741] <= 32'b00000000000000000000000000000000;
REG[742] <= 32'b00000000000000000000000000001010;
REG[743] <= 32'b00001011000000000000000100001101;
REG[744] <= 32'b00000000000000000000000000000000;
REG[745] <= 32'b00000000000000000000000000000000;
REG[746] <= 32'b00000000000000000000000000000000;
REG[747] <= 32'b00000000000000000001011100000000;
REG[748] <= 32'b00000000000000000000000000000000;
REG[749] <= 32'b00000000000000000001101000000011;
REG[750] <= 32'b00000000000000000000000000000000;
REG[751] <= 32'b00000000000000000000000000000000;
REG[752] <= 32'b00000000000000000001011100000000;
REG[753] <= 32'b00000000000000000000000000000000;
REG[754] <= 32'b00000000000000000000000000000000;
REG[755] <= 32'b00000000000000000001100100000000;
REG[756] <= 32'b00000000000000000000000000000000;
REG[757] <= 32'b00000000000000000000000000000000;
REG[758] <= 32'b00000000000000000000000000000000;
REG[759] <= 32'b00000000000000000000000000000000;
REG[760] <= 32'b00000000000000000000000000000000;
REG[761] <= 32'b00000000000000000000000000000000;
REG[762] <= 32'b00000000000000000000000000000000;
REG[763] <= 32'b00000000000000000000000000000000;
REG[764] <= 32'b00000000000000000000000000011001;
REG[765] <= 32'b00000000000000000000000000000000;
REG[766] <= 32'b00000000000001000010010100101010;
REG[767] <= 32'b00000000000000000000000000101010;
REG[768] <= 32'b00000000000000000000000000000000;
REG[769] <= 32'b00000000000000000000000000000000;
REG[770] <= 32'b00000000000000000000000000000000;
REG[771] <= 32'b00000000000010100000000000000000;
REG[772] <= 32'b00000000000000000000000000000000;
REG[773] <= 32'b00000000000000000000000000000000;
REG[774] <= 32'b00000000000000000000000000000000;
REG[775] <= 32'b00000000000000000000000000000000;
REG[776] <= 32'b00000000000000000000000000000000;
REG[777] <= 32'b00000000000011110000000000000000;
REG[778] <= 32'b00000000000000010000000000000000;
REG[779] <= 32'b00000000000000000000000000000000;
REG[780] <= 32'b00000000000000000000000000000000;
REG[781] <= 32'b00000000000000000000000000000000;
REG[782] <= 32'b00000000000000000000000000000000;
REG[783] <= 32'b00000000000000000000000000000000;
REG[784] <= 32'b00000000000000000000000000010010;
REG[785] <= 32'b00011011000001110001011100000101;
REG[786] <= 32'b00000000000000000000000000000000;
REG[787] <= 32'b00000000000000000001010000010100;
REG[788] <= 32'b00000000000000000001111100010000;
REG[789] <= 32'b00000000000000000000000000000000;
REG[790] <= 32'b00000000000000000001010000010010;
REG[791] <= 32'b00000000000000110010001000001110;
REG[792] <= 32'b00000000000000000000000000000000;
REG[793] <= 32'b00000000000000000000000000000000;
REG[794] <= 32'b00000000000000000000000000000000;
REG[795] <= 32'b00000000000000000000000000000000;
REG[796] <= 32'b00100010001001010000000000000000;
REG[797] <= 32'b00010010000000000000000000001110;
REG[798] <= 32'b00000000000101010000000000000000;
REG[799] <= 32'b00000000000000000000000000001011;
REG[800] <= 32'b00000101000000000000000000000000;
REG[801] <= 32'b00000000001010100000000000000000;
REG[802] <= 32'b00001100000011100000000000001100;
REG[803] <= 32'b00010000000000000000000000000000;
REG[804] <= 32'b00000000000000000000000000000000;
REG[805] <= 32'b00000000000000000000000000000000;
REG[806] <= 32'b00000000000000000000000000000000;
REG[807] <= 32'b00000000000000000000000000110000;
REG[808] <= 32'b00101101001011000011001000000110;
REG[809] <= 32'b00000000000000000000000000000000;
REG[810] <= 32'b00000000000000000000000000000000;
REG[811] <= 32'b00000000000000000000000000000011;
REG[812] <= 32'b00101000000000000000000000000000;
REG[813] <= 32'b00000000000001100000100000000000;
REG[814] <= 32'b00000000000001110001101100100100;
REG[815] <= 32'b00101001000000000000000000000000;
REG[816] <= 32'b00000000000000000000000000000000;
REG[817] <= 32'b00000000000000000000000000000000;
REG[818] <= 32'b00000000000000000000000000000000;
REG[819] <= 32'b00000000000001110000000000000000;
REG[820] <= 32'b00000000000000000000000000000000;
REG[821] <= 32'b00000000000000000000000000010100;
REG[822] <= 32'b00000000000000000000000000000000;
REG[823] <= 32'b00000000000000000000000000000000;
REG[824] <= 32'b00000010000000000000000000100110;
REG[825] <= 32'b00000000000010000000000000000000;
REG[826] <= 32'b00100110000000000000000000001001;
REG[827] <= 32'b00001001000000000000000000000000;
REG[828] <= 32'b00000000000000000000000000000000;
REG[829] <= 32'b00000000000000000000000000000000;
REG[830] <= 32'b00000000000000000000000000000000;
REG[831] <= 32'b00000000000000100001000100000000;
REG[832] <= 32'b00000000000000000001110100011110;
REG[833] <= 32'b00000011000000110000000000000000;
REG[834] <= 32'b00000000000000000000000000000000;
REG[835] <= 32'b00000000000000000011001000000000;
REG[836] <= 32'b00000000000111000000000100000111;
REG[837] <= 32'b00000000000000110000110000000000;
REG[838] <= 32'b00000000000000000011001000011001;
REG[839] <= 32'b00000100000000000001000000010101;
REG[840] <= 32'b00000000000000000000000000000000;
REG[841] <= 32'b00000000000000000000000000000000;
REG[842] <= 32'b00000000000000000000000000000000;
REG[843] <= 32'b00000000000000000000101000000000;
REG[844] <= 32'b00000000000000000000000000010010;
REG[845] <= 32'b00000101000000000000000000000000;
REG[846] <= 32'b00000000000000000000000000000000;
REG[847] <= 32'b00000000000000000000000000010101;
REG[848] <= 32'b00000000000000000000000000000000;
REG[849] <= 32'b00000000000000000000000000000000;
REG[850] <= 32'b00000100000000000000000000011000;
REG[851] <= 32'b00000000000000000000011000000000;
REG[852] <= 32'b00000000000000000000000000000000;
REG[853] <= 32'b00000000000000000000000000000000;
REG[854] <= 32'b00000000000000000000000000000000;
REG[855] <= 32'b00010111000000110000000000000000;
REG[856] <= 32'b00000000000000000000010000000000;
REG[857] <= 32'b00000000000000000000000000000000;
REG[858] <= 32'b00010100000010100000000000000000;
REG[859] <= 32'b00000000000000000000000000000000;
REG[860] <= 32'b00000000000000000000110100001010;
REG[861] <= 32'b00001110000011110000000000000000;
REG[862] <= 32'b00000000000000000000000000000000;
REG[863] <= 32'b00000000000000000000011000001111;
REG[864] <= 32'b00000000000000000000000000000000;
REG[865] <= 32'b00000000000000000000000000000000;
REG[866] <= 32'b00000000000000000000000000000000;
REG[867] <= 32'b00000000000000000000000000000000;
REG[868] <= 32'b00000000000000000000000000000000;
REG[869] <= 32'b00000000000000000000000000000010;
REG[870] <= 32'b00000000000000000000000000000000;
REG[871] <= 32'b00000000000000000000000000000000;
REG[872] <= 32'b00000000000000000000000000000000;
REG[873] <= 32'b00000000000000000000000000000000;
REG[874] <= 32'b00000000000000000000000000000000;
REG[875] <= 32'b00000000000000000000000000000000;
REG[876] <= 32'b00000000000000000000000000000000;
REG[877] <= 32'b00000000000000000000000000000000;
REG[878] <= 32'b00000000000000000000000000000000;
REG[879] <= 32'b00000000000000000000000000000011;
REG[880] <= 32'b00000000000000000000000000000000;
REG[881] <= 32'b00000000000001000000000000000000;
REG[882] <= 32'b00000000000000000000101000000000;
REG[883] <= 32'b00010111000011100000000000000000;
REG[884] <= 32'b00000000000000000000000000000000;
REG[885] <= 32'b00000000000000000000000000000000;
REG[886] <= 32'b00000000000000000000000000000000;
REG[887] <= 32'b00000000000000000000000000000000;
REG[888] <= 32'b00000000000000000000000000000000;
REG[889] <= 32'b00000000000000000000000000000000;
REG[890] <= 32'b00000000000000000000000000000000;
REG[891] <= 32'b00000000001101010000110100000000;
REG[892] <= 32'b00000000000000000000000000001101;
REG[893] <= 32'b00000000000000000000000000000001;
REG[894] <= 32'b00000000000111000000000000000000;
REG[895] <= 32'b00000000000000000000000000100100;
REG[896] <= 32'b00011010000000000000000000010101;
REG[897] <= 32'b00000000001000110000000000000000;
REG[898] <= 32'b00001001000001000000000000000110;
REG[899] <= 32'b00000000000000000000000000000000;
REG[900] <= 32'b00000000000000000000000000000000;
REG[901] <= 32'b00000000000000000000000000000000;
REG[902] <= 32'b00000000000000000000000000000000;
REG[903] <= 32'b00010100000101110001110000000000;
REG[904] <= 32'b00000000000000000000000000000011;
REG[905] <= 32'b00000000000000100000000000000000;
REG[906] <= 32'b00000000000000000000000000000000;
REG[907] <= 32'b00001011000011110000000000000000;
REG[908] <= 32'b00000100001000000000011100000000;
REG[909] <= 32'b00000001000110100000000000001101;
REG[910] <= 32'b00001001000001100000000000000000;
REG[911] <= 32'b00000101000000000000000000000000;
REG[912] <= 32'b00000000000000000000000000000000;
REG[913] <= 32'b00000000000000000000000000000000;
REG[914] <= 32'b00000000000000000000000000000000;
REG[915] <= 32'b00000000000011110001111000000000;
REG[916] <= 32'b00001110000000000000000000100000;
REG[917] <= 32'b01001000000000000000000000010000;
REG[918] <= 32'b00000000000000110000000000000000;
REG[919] <= 32'b00000000000000000000000000000000;
REG[920] <= 32'b00011010000000000000000000000000;
REG[921] <= 32'b00000000000000000000000000000000;
REG[922] <= 32'b00010100000000000000000000000000;
REG[923] <= 32'b00000001000000000000000000000000;
REG[924] <= 32'b00000000000000000000000000000000;
REG[925] <= 32'b00000000000000000000000000000000;
REG[926] <= 32'b00000000000000000000000000000000;
REG[927] <= 32'b00011111000000000000000000000000;
REG[928] <= 32'b00000000000000000010101000011010;
REG[929] <= 32'b00101100001011010000111000000000;
REG[930] <= 32'b00011001000100000000000000000000;
REG[931] <= 32'b00000000000000000000000100000000;
REG[932] <= 32'b00000000000110010000011100000000;
REG[933] <= 32'b00000000000000000000000000000000;
REG[934] <= 32'b00000000000000000000000000000000;
REG[935] <= 32'b00000000001011100001110000000000;
REG[936] <= 32'b00000000000000000000000000000000;
REG[937] <= 32'b00000000000000000000000000000000;
REG[938] <= 32'b00000000000000000000000000000000;
REG[939] <= 32'b00000000000000000000000000000000;
REG[940] <= 32'b00001110000011110000000000000000;
REG[941] <= 32'b00000000000000000000000000000000;
REG[942] <= 32'b00000000000010000000000000000000;
REG[943] <= 32'b00000000000000000000000000000000;
REG[944] <= 32'b00000000000000000000101100000000;
REG[945] <= 32'b00000000000110000000000000000000;
REG[946] <= 32'b00000000000000000000000000001100;
REG[947] <= 32'b00000000000000000000010100000000;
REG[948] <= 32'b00000000000000000000000000000000;
REG[949] <= 32'b00000000000000000000000000000000;
REG[950] <= 32'b00000000000000000000000000000000;
REG[951] <= 32'b00001011000111110000000000000000;
REG[952] <= 32'b00000000000000000001001000001101;
REG[953] <= 32'b00000000000000000000000000000000;
REG[954] <= 32'b00000000001000110001010000011000;
REG[955] <= 32'b00001000000000000000000000011110;
REG[956] <= 32'b00000000000000000000000000000000;
REG[957] <= 32'b00000000000111110000111000010111;
REG[958] <= 32'b00000000000000000000000000001100;
REG[959] <= 32'b00000011000000000000000000000000;
REG[960] <= 32'b00000000000000000000000000000000;
REG[961] <= 32'b00000000000000000000000000000000;
REG[962] <= 32'b00000000000000000000000000000000;
REG[963] <= 32'b00000000000010000011100000000000;
REG[964] <= 32'b00100011000101000000000000000000;
REG[965] <= 32'b00000000000000000000000000000000;
REG[966] <= 32'b00000000000000000011010100000000;
REG[967] <= 32'b00100101000000000000000000000000;
REG[968] <= 32'b00000000000000000000000000000000;
REG[969] <= 32'b00000000000000000000000000000000;
REG[970] <= 32'b00101110000000000000000000000000;
REG[971] <= 32'b00000000000000000010010100000000;
REG[972] <= 32'b00000000000000000000000000000000;
REG[973] <= 32'b00000000000000000000000000000000;
REG[974] <= 32'b00000000000000000000000000000000;
REG[975] <= 32'b00000000000000000000000000100010;
REG[976] <= 32'b00101011001100000000000000000000;
REG[977] <= 32'b00000000000000000000000000000000;
REG[978] <= 32'b00100111000000000000000000000000;
REG[979] <= 32'b00011100000111000000000000000000;
REG[980] <= 32'b00000000000000000000000000000000;
REG[981] <= 32'b00000000000000000000000000000000;
REG[982] <= 32'b00001110000011000000000000000000;
REG[983] <= 32'b00000000000000000000000000000000;
REG[984] <= 32'b00000000000000000000000000000000;
REG[985] <= 32'b00000000000000000000000000000000;
REG[986] <= 32'b00000000000000000000000000000000;
REG[987] <= 32'b00000000000111010011010100000000;
REG[988] <= 32'b00000110000111000000000000000000;
REG[989] <= 32'b00010011000000000000000100010110;
REG[990] <= 32'b00000000000000000000010100000000;
REG[991] <= 32'b00001011000001000000000000000101;
REG[992] <= 32'b00001110000000000000000000011011;
REG[993] <= 32'b00000000000000000000000000000000;
REG[994] <= 32'b00010100000101010000000000000000;
REG[995] <= 32'b00000000000000000000000000011100;
REG[996] <= 32'b00000000000000000000000000000000;
REG[997] <= 32'b00000000000000000000000000000000;
REG[998] <= 32'b00000000000000000000000000000000;
REG[999] <= 32'b00000000000000000001111000100100;
REG[1000] <= 32'b00000110000001100000000000000000;
REG[1001] <= 32'b00011000000000000000000000000000;
REG[1002] <= 32'b00000000000010100000110100001100;
REG[1003] <= 32'b00000110000100100001010000000000;
REG[1004] <= 32'b00000000000000000000000000000000;
REG[1005] <= 32'b00000000000000000000101000010010;
REG[1006] <= 32'b00000000000000000001100000000000;
REG[1007] <= 32'b00000000000010000000000000000000;
REG[1008] <= 32'b00000000000000000000000000000000;
REG[1009] <= 32'b00000000000000000000000000000000;
REG[1010] <= 32'b00000000000000000000000000000000;
REG[1011] <= 32'b00000000000000000000000000000000;
REG[1012] <= 32'b00000000000000000000000000001010;
REG[1013] <= 32'b00100101000000000000111100000011;
REG[1014] <= 32'b00000000000000000000000000000000;
REG[1015] <= 32'b00100111000000000000000000000000;
REG[1016] <= 32'b00000000000000000001100100000000;
REG[1017] <= 32'b00000000000000000000000000000000;
REG[1018] <= 32'b00011111000000000000000000000000;
REG[1019] <= 32'b00000000000000000010110100000000;
REG[1020] <= 32'b00000000000000000000000000000000;
REG[1021] <= 32'b00000000000000000000000000000000;
REG[1022] <= 32'b00000000000000000000000000000000;
REG[1023] <= 32'b00000000000000000010010100000000;
REG[1024] <= 32'b00000111000011000010101000001011;
REG[1025] <= 32'b00010101000000000000000000011000;
REG[1026] <= 32'b00000000000000000001011000000000;
REG[1027] <= 32'b01000100010101010000000000000000;
REG[1028] <= 32'b00010100000000000000000000101100;
REG[1029] <= 32'b00000000000000000000000000000000;
REG[1030] <= 32'b00101110010010010000000000001110;
REG[1031] <= 32'b00010100000000000000000000000000;
REG[1032] <= 32'b00000000000000000000000000000000;
REG[1033] <= 32'b00000000000000000000000000000000;
REG[1034] <= 32'b00000000000000000000000000000000;
REG[1035] <= 32'b00000000000000000000000000000000;
REG[1036] <= 32'b00000000000000000000000000000000;
REG[1037] <= 32'b00011010000000000000000000000000;
REG[1038] <= 32'b00000000000000000000000000000000;
REG[1039] <= 32'b00010010000000000000000000000000;
REG[1040] <= 32'b00100001000000000000000000000000;
REG[1041] <= 32'b00000000000000000000000000000000;
REG[1042] <= 32'b00000000000000000000000000000000;
REG[1043] <= 32'b00000000000000000000000000000000;
REG[1044] <= 32'b00000000000000000000000000000000;
REG[1045] <= 32'b00000000000000000000000000000000;
REG[1046] <= 32'b00000000000000000000000000000000;
REG[1047] <= 32'b00010010000011000000000000000000;
REG[1048] <= 32'b00000000000000000000110100000000;
REG[1049] <= 32'b00000000000000000000001100000000;
REG[1050] <= 32'b00000000001101000001001100000000;
REG[1051] <= 32'b00000000000000000011001100000000;
REG[1052] <= 32'b00000000000000000010111100001001;
REG[1053] <= 32'b00000000000100100000000100000000;
REG[1054] <= 32'b00000000000000000001111000001111;
REG[1055] <= 32'b00000000000001010010011100010000;
REG[1056] <= 32'b00000000000000000000000000000000;
REG[1057] <= 32'b00000000000000000000000000000000;
REG[1058] <= 32'b00000000000000000000000000000000;
REG[1059] <= 32'b00000000000001010000001100000000;
REG[1060] <= 32'b00000000000011110000000000000000;
REG[1061] <= 32'b00000000000000000010111100010011;
REG[1062] <= 32'b00000000001010000011001000000000;
REG[1063] <= 32'b00000000000000000000000000000011;
REG[1064] <= 32'b00000000000000000010101100010011;
REG[1065] <= 32'b00000000001110100100111100000000;
REG[1066] <= 32'b00000000000000000000000000000000;
REG[1067] <= 32'b00000000000000000000101000000010;
REG[1068] <= 32'b00000000000000000000000000000000;
REG[1069] <= 32'b00000000000000000000000000000000;
REG[1070] <= 32'b00000000000000000000000000000000;
REG[1071] <= 32'b00001010000111000010000000000000;
REG[1072] <= 32'b00000000000000000000000000000000;
REG[1073] <= 32'b00000000000111010010100000101000;
REG[1074] <= 32'b00100001000100100001111000000000;
REG[1075] <= 32'b00000000000000000000000000000000;
REG[1076] <= 32'b00000000000010010000000000000000;
REG[1077] <= 32'b00011101000001010000110000000000;
REG[1078] <= 32'b00000000000000000000000000000000;
REG[1079] <= 32'b00000000000101100000000000000000;
REG[1080] <= 32'b00000000000000000000000000000000;
REG[1081] <= 32'b00000000000000000000000000000000;
REG[1082] <= 32'b00000000000000000000000000000000;
REG[1083] <= 32'b00000000000010010001011000000000;
REG[1084] <= 32'b00000000000010010000000000000110;
REG[1085] <= 32'b00011011000000000000000000000000;
REG[1086] <= 32'b00000000001100010001001000000000;
REG[1087] <= 32'b00000011000000000000000000000000;
REG[1088] <= 32'b00000000000000000000000000000000;
REG[1089] <= 32'b00000000000110010001111100000000;
REG[1090] <= 32'b00010100000000000000000000000000;
REG[1091] <= 32'b00000000000000000000000000000000;
REG[1092] <= 32'b00000000000000000000000000000000;
REG[1093] <= 32'b00000000000000000000000000000000;
REG[1094] <= 32'b00000000000000000000000000000000;
REG[1095] <= 32'b00010000000000000000000000011110;
REG[1096] <= 32'b00010011000000000001100100000000;
REG[1097] <= 32'b00000000000000000000000000000000;
REG[1098] <= 32'b00000000000000000000001100000000;
REG[1099] <= 32'b00011010000010100000000000000000;
REG[1100] <= 32'b00000000000000000000000000000000;
REG[1101] <= 32'b00010011000000000000000000000000;
REG[1102] <= 32'b00010110000011010000000000001001;
REG[1103] <= 32'b00000000000000000000000000000000;
REG[1104] <= 32'b00000000000000000000000000000000;
REG[1105] <= 32'b00000000000000000000000000000000;
REG[1106] <= 32'b00000000000000000000000000000000;
REG[1107] <= 32'b00000000000000000000000000000000;
REG[1108] <= 32'b00000000000101100000000000110010;
REG[1109] <= 32'b00000000000000000100101100110011;
REG[1110] <= 32'b00000000000000000000000000000000;
REG[1111] <= 32'b00000000000000000000000000010011;
REG[1112] <= 32'b00000001000000000000100100000000;
REG[1113] <= 32'b00000000000000000000000000000000;
REG[1114] <= 32'b00001001000000000000000000000000;
REG[1115] <= 32'b00000000000000000001010100000000;
REG[1116] <= 32'b00000000000000000000000000000000;
REG[1117] <= 32'b00000000000000000000000000000000;
REG[1118] <= 32'b00000000000000000000000000000000;
REG[1119] <= 32'b00000000000000000000000000001110;
REG[1120] <= 32'b00000000000000000000000000000000;
REG[1121] <= 32'b00000000010101110101110101010000;
REG[1122] <= 32'b00001110000000000000000000000000;
REG[1123] <= 32'b00000000000000000000000000000000;
REG[1124] <= 32'b00000000000000000000000000000000;
REG[1125] <= 32'b00001011000100000000000000000000;
REG[1126] <= 32'b00000000000000000000000000000000;
REG[1127] <= 32'b00000000000000000000100000010101;
REG[1128] <= 32'b00000000000000000000000000000000;
REG[1129] <= 32'b00000000000000000000000000000000;
REG[1130] <= 32'b00000000000000000000000000000000;
REG[1131] <= 32'b00000000000101000000110000000000;
REG[1132] <= 32'b00000000000000000000000000000000;
REG[1133] <= 32'b00000000000000000000111000011100;
REG[1134] <= 32'b00000000000000000000000000000000;
REG[1135] <= 32'b00000000000000000000000000000000;
REG[1136] <= 32'b00000000000000000000000000000000;
REG[1137] <= 32'b00000000000000000000000000000000;
REG[1138] <= 32'b00000000000000000000000000000000;
REG[1139] <= 32'b00000000000000000000000000000000;
REG[1140] <= 32'b00000000000000000000000000000000;
REG[1141] <= 32'b00000000000000000000000000000000;
REG[1142] <= 32'b00000000000000000000000000000000;
REG[1143] <= 32'b00000000000011010000101000000000;
REG[1144] <= 32'b00000000000000000000000000000000;
REG[1145] <= 32'b00000000000000110000000000000000;
REG[1146] <= 32'b00000000000000000000000000000000;
REG[1147] <= 32'b00000000000000000000000000000000;
REG[1148] <= 32'b00000000000000000000000000000000;
REG[1149] <= 32'b00000000000000000000001100000000;
REG[1150] <= 32'b00000000000000000000000000000000;
REG[1151] <= 32'b00000000000000000000000000000000;







////////////////////////////////////////////////////
//// FILTER
////////////////////////////////////////////////////




REG[2040] <= 32'b0;
REG[2041] <= 32'b0;
REG[2042] <= 32'b0;
REG[2043] <= 32'b0;
REG[2044] <= 32'b0;
REG[2045] <= 32'b0;
REG[2046] <= 32'b0;
REG[2047] <= 32'b0;
REG[2048] <= 32'b0;
REG[2049] <= 32'b0;
REG[2050] <= 32'b0;
REG[2051] <= 32'b0;
REG[2052] <= 32'b0;
REG[2053] <= 32'b0;
REG[2054] <= 32'b0;
REG[2055] <= 32'b0;
REG[2056] <= 32'b0;
REG[2057] <= 32'b0;
REG[2058] <= 32'b0;
REG[2059] <= 32'b0;
REG[2060] <= 32'b0;
REG[2061] <= 32'b0;
REG[2062] <= 32'b0;
REG[2063] <= 32'b0;
REG[2064] <= 32'b1111_1100_0001_1001_0000_0001_0000_0000;
REG[2065] <= 32'b00000011000011010000010100101101;
REG[2066] <= 32'b00001110111110110000000000000001;
REG[2067] <= 32'b11111100000101010000000011110001;
REG[2068] <= 32'b11110100111110001111100100000010;
REG[2069] <= 32'b00000000111111111111000111111011;
REG[2070] <= 32'b00000111000010111111110000001001;
REG[2071] <= 32'b11110100111111010000001000000100;
REG[2072] <= 32'b00000101000000011111000111111001;
REG[2073] <= 32'b11101010000010100000010111111001;
REG[2074] <= 32'b11111001111111101110100100011000;
REG[2075] <= 32'b00010101000001010000000111111001;
REG[2076] <= 32'b11101010111110011111110111111010;
REG[2077] <= 32'b00000101000000011111110011111011;
REG[2078] <= 32'b11110011111111110000010011111101;
REG[2079] <= 32'b11101101111011111111001000000101;
REG[2080] <= 32'b00000001111111111110111111101100;
REG[2081] <= 32'b00000000111101110000000111111111;
REG[2082] <= 32'b00000010000001010000110000000110;
REG[2083] <= 32'b00000100000010100000010100000000;
REG[2084] <= 32'b00001000111110110000110000011011;
REG[2085] <= 32'b00010010000001110000111111111111;
REG[2086] <= 32'b00001000001000101111101011110010;
REG[2087] <= 32'b11110111111101100000001111111110;
REG[2088] <= 32'b11110100111100111111011111101100;
REG[2089] <= 32'b11111100000001101110111011101110;
REG[2090] <= 32'b11101010111100011111110100000010;
REG[2091] <= 32'b11111111000001010000101011110111;
REG[2092] <= 32'b00000011000011011111010011111100;
REG[2093] <= 32'b00000101111101111111110100000000;
REG[2094] <= 32'b11110111111110011111111111110111;
REG[2095] <= 32'b11111000111111001110111111101101;
REG[2096] <= 32'b11110000111111000001001000010100;
REG[2097] <= 32'b00000000000001011111110111110011;
REG[2098] <= 32'b00000101000101001111110100000001;
REG[2099] <= 32'b00000101111110010000010100001011;
REG[2100] <= 32'b00000100111100111111100111111000;
REG[2101] <= 32'b11110101111110000000011011110100;
REG[2102] <= 32'b11111001111111101111010011111100;
REG[2103] <= 32'b11111010111101010000000111111110;
REG[2104] <= 32'b11110101000001001111001011101100;
REG[2105] <= 32'b00001001111101101111010100000000;
REG[2106] <= 32'b11111000111110110000011111110100;
REG[2107] <= 32'b11111001000000111111000011111110;
REG[2108] <= 32'b00001001111100111111010111110111;
REG[2109] <= 32'b11110101111110010000011100000010;
REG[2110] <= 32'b11111000111101001110101011101110;
REG[2111] <= 32'b11111011000000111111011011101110;
REG[2112] <= 32'b11101110111101101111100100000101;
REG[2113] <= 32'b11110100111101011111011100000000;
REG[2114] <= 32'b11111001111110000000010100001100;
REG[2115] <= 32'b00001001000100100000001111101110;
REG[2116] <= 32'b00000111000011100000110100010011;
REG[2117] <= 32'b11110010111101100000011100000111;
REG[2118] <= 32'b11101111110111011111011011101110;
REG[2119] <= 32'b00001010000100101111010011100011;
REG[2120] <= 32'b11110111111101110001001000011001;
REG[2121] <= 32'b11101101111011010000001011110100;
REG[2122] <= 32'b11111011000000011111100100010011;
REG[2123] <= 32'b00011000111101011111100100000001;
REG[2124] <= 32'b00000010000111110001111011110100;
REG[2125] <= 32'b11110100111110001111000000000010;
REG[2126] <= 32'b11111011111101001111000011110101;
REG[2127] <= 32'b00000101000011000001000100001000;
REG[2128] <= 32'b00001001000100110000111000010100;
REG[2129] <= 32'b00001100111111111111111100000001;
REG[2130] <= 32'b00010100000101100001010100000010;
REG[2131] <= 32'b11111010111110001110110111110100;
REG[2132] <= 32'b11110101000001000001000100000111;
REG[2133] <= 32'b11101110111100111111100000010110;
REG[2134] <= 32'b00110011001010101110100011101110;
REG[2135] <= 32'b11110100000010010001001100001000;
REG[2136] <= 32'b11110011111000111111011011111001;
REG[2137] <= 32'b11110110111110111111011011101011;
REG[2138] <= 32'b11111010111111001111011111111010;
REG[2139] <= 32'b00000000111100001111101100000000;
REG[2140] <= 32'b11111010000001001111001100011101;
REG[2141] <= 32'b11111110000000010000110100010001;
REG[2142] <= 32'b00000011000111001111000111111011;
REG[2143] <= 32'b00000010000001000010010000011100;
REG[2144] <= 32'b11100100000000100000011100001001;
REG[2145] <= 32'b11110011000000100001111111110011;
REG[2146] <= 32'b11110110111101101110100011101011;
REG[2147] <= 32'b00000010111011101111000011111011;
REG[2148] <= 32'b11101100111101010000010011110111;
REG[2149] <= 32'b11111100000001000000011011101110;
REG[2150] <= 32'b11101110000010001111110011111111;
REG[2151] <= 32'b00000011111110111111111000000011;
REG[2152] <= 32'b11111011111110101111101011111010;
REG[2153] <= 32'b00000110000000011111111011111111;
REG[2154] <= 32'b00010000111101111110111111110111;
REG[2155] <= 32'b11110001111100100000010011110001;
REG[2156] <= 32'b11101101111110011111001011110110;
REG[2157] <= 32'b11101110111100011111011000000100;
REG[2158] <= 32'b11111110111110011111100000010001;
REG[2159] <= 32'b00010101000101100000110111111011;
REG[2160] <= 32'b11110110000101100000100000010001;
REG[2161] <= 32'b00001101111111100000011011111110;
REG[2162] <= 32'b11101001000101010000101100000011;
REG[2163] <= 32'b00010001000010000000101000001010;
REG[2164] <= 32'b00001101000011000001000000001010;
REG[2165] <= 32'b00001010111101010000010000000000;
REG[2166] <= 32'b11110111111111100000101100001011;
REG[2167] <= 32'b00001000111100110000100000000111;
REG[2168] <= 32'b11111111111101000000010100001001;
REG[2169] <= 32'b00000001000100001111111000000001;
REG[2170] <= 32'b00000111000010010000100100011010;
REG[2171] <= 32'b00001010000011000001100100010110;
REG[2172] <= 32'b11101000111101101111010111110010;
REG[2173] <= 32'b11101110000010011110011011101111;
REG[2174] <= 32'b00000010111100001111000100000110;
REG[2175] <= 32'b11101111000001010000001111101011;
REG[2176] <= 32'b11101111000000000001000000000101;
REG[2177] <= 32'b00000000111110010000001111111111;
REG[2178] <= 32'b11111100111110010000000111110110;
REG[2179] <= 32'b00000010000001111111100111110101;
REG[2180] <= 32'b00000000111100011111110000000011;
REG[2181] <= 32'b00000011000010010010011011110100;
REG[2182] <= 32'b00000001111011000000101000001001;
REG[2183] <= 32'b00010111111101100000010111101101;
REG[2184] <= 32'b11111111000000110000100011110010;
REG[2185] <= 32'b00000001111010011111001000100110;
REG[2186] <= 32'b00001010000000000000000000000100;
REG[2187] <= 32'b00010010001100101111110100000011;
REG[2188] <= 32'b00000001000000000001010100010011;
REG[2189] <= 32'b11110110000011000000101000000000;
REG[2190] <= 32'b11111100000001010000110011110110;
REG[2191] <= 32'b11110110000001011111100100000000;
REG[2192] <= 32'b00000010111110111111110111111100;
REG[2193] <= 32'b11111101111111101111110000000000;
REG[2194] <= 32'b00000100000000000000011000000000;
REG[2195] <= 32'b11101110000000001111111011111101;
REG[2196] <= 32'b11110110111110011111000011110011;
REG[2197] <= 32'b11110100111110001110110011111011;
REG[2198] <= 32'b11110101111100111111001111111010;
REG[2199] <= 32'b11111001111111101111111111111000;
REG[2200] <= 32'b00001000000100011111111100000011;
REG[2201] <= 32'b00000111111101000000010000000101;
REG[2202] <= 32'b00000010000001010000100111110111;
REG[2203] <= 32'b00000100111110111111100011101100;
REG[2204] <= 32'b11111001111101101111000011110101;
REG[2205] <= 32'b11101100111101010000000000000000;
REG[2206] <= 32'b11111010000000001110110011110111;
REG[2207] <= 32'b11111010000001101111111000000110;
REG[2208] <= 32'b11110011111111010000001100010001;
REG[2209] <= 32'b00001110000011110000010000001010;
REG[2210] <= 32'b11111011111111110000000111111010;
REG[2211] <= 32'b00001111000101111111101011111101;
REG[2212] <= 32'b11111111111110011111110011111100;
REG[2213] <= 32'b00000110000000111111110011110011;
REG[2214] <= 32'b11111100111101100000000000101011;
REG[2215] <= 32'b00000101111101101111111111111000;
REG[2216] <= 32'b00000001001011000001100111110111;
REG[2217] <= 32'b11100000000000101111110011101111;
REG[2218] <= 32'b11101100000000011111110011101001;
REG[2219] <= 32'b11101111111010101110111100001110;
REG[2220] <= 32'b00000110111110000000100011111011;
REG[2221] <= 32'b00000011000100011110111111111010;
REG[2222] <= 32'b00000111111101110000100100010100;
REG[2223] <= 32'b11101001111011101111111000010110;
REG[2224] <= 32'b11110111000010101111001111110111;
REG[2225] <= 32'b00000000111011101111100000010000;
REG[2226] <= 32'b00000000000011110000110011110110;
REG[2227] <= 32'b11111011111111010000000011111111;
REG[2228] <= 32'b11111001111111110001000100000000;
REG[2229] <= 32'b11111110000000001111101100000111;
REG[2230] <= 32'b00000111111110101111111011111100;
REG[2231] <= 32'b11111010111111001111100011111111;
REG[2232] <= 32'b11111001111101001110111111110011;
REG[2233] <= 32'b11110111000000001111010111101111;
REG[2234] <= 32'b11110100111100111111100111111010;
REG[2235] <= 32'b11110101111101100000100011111001;
REG[2236] <= 32'b00000011000011011111000000000000;
REG[2237] <= 32'b00001110111100101111101111110100;
REG[2238] <= 32'b11101011111101100000100011110111;
REG[2239] <= 32'b11111011111101111111110111110100;
REG[2240] <= 32'b11111011000010010010010100011111;
REG[2241] <= 32'b11111101111101001111011000010010;
REG[2242] <= 32'b00010001000100100000001111110101;
REG[2243] <= 32'b11110111000001100000000000000011;
REG[2244] <= 32'b11100010111010110000110000010000;
REG[2245] <= 32'b00000111111110111111100000010010;
REG[2246] <= 32'b11111000111110101110110111110000;
REG[2247] <= 32'b00010000000010101110011000000100;
REG[2248] <= 32'b11111100111111010000001100000000;
REG[2249] <= 32'b00010011111111101111011111110010;
REG[2250] <= 32'b00000010111101011111110100101101;
REG[2251] <= 32'b00100110111101000000001000000111;
REG[2252] <= 32'b00000101111100111111110011110100;
REG[2253] <= 32'b11111010111110010000001000000001;
REG[2254] <= 32'b11111010000000011111101100000000;
REG[2255] <= 32'b11111110111111011111000111110101;
REG[2256] <= 32'b00001110000101010000110100001000;
REG[2257] <= 32'b00000000111110101111010111111101;
REG[2258] <= 32'b00001010111101011110111111111100;
REG[2259] <= 32'b11111111111011110000001000010010;
REG[2260] <= 32'b00000110111100010000100100000110;
REG[2261] <= 32'b00010101000011010000101011111101;
REG[2262] <= 32'b11111100111101011111001111111111;
REG[2263] <= 32'b00000111000100010001001111111111;
REG[2264] <= 32'b11111101111110000001001000100011;
REG[2265] <= 32'b11111000111111110000011011110101;
REG[2266] <= 32'b00000111111111101111011100001001;
REG[2267] <= 32'b11110101111110011111111111111101;
REG[2268] <= 32'b11101111000000011111100111110110;
REG[2269] <= 32'b11111000000001000000011000000100;
REG[2270] <= 32'b11111010111101101111010011111001;
REG[2271] <= 32'b11110000111101101111000011101100;
REG[2272] <= 32'b11101011111011011110110111101001;
REG[2273] <= 32'b11101111111011111111010011110001;
REG[2274] <= 32'b11100010111011101110110011110001;
REG[2275] <= 32'b11110101111101111110111111111111;
REG[2276] <= 32'b00000011111110101111100011110001;
REG[2277] <= 32'b11111111000101100000111011101101;
REG[2278] <= 32'b11101011111101111111010011111101;
REG[2279] <= 32'b00000100111010111110111011110010;
REG[2280] <= 32'b00001010000100010001000100001100;
REG[2281] <= 32'b00000101111101110001000100011010;
REG[2282] <= 32'b11111101000010011111001011100110;
REG[2283] <= 32'b00001100000001010000110111111101;
REG[2284] <= 32'b11110100111111101111110011101111;
REG[2285] <= 32'b11110111000010110001010000000000;
REG[2286] <= 32'b11110011111001111110110000011000;
REG[2287] <= 32'b00010110111110100000000111110111;
REG[2288] <= 32'b00000010000011011110111111101101;
REG[2289] <= 32'b11111100111101010000000011111111;
REG[2290] <= 32'b11111100111101010001001000001000;
REG[2291] <= 32'b11110100000000000000000011101110;
REG[2292] <= 32'b00010110000011100000010000010001;
REG[2293] <= 32'b00001110111100010000000000000000;
REG[2294] <= 32'b11110101111110001111111000000001;
REG[2295] <= 32'b11111010111110011111000000001010;
REG[2296] <= 32'b11110000111111011111011011110010;
REG[2297] <= 32'b11110011111101001111001011111000;
REG[2298] <= 32'b11101101111100001111001111111010;
REG[2299] <= 32'b00000001000000101111111000001001;
REG[2300] <= 32'b00001001000000110001100000010110;
REG[2301] <= 32'b00000010000110100001010000001001;
REG[2302] <= 32'b00001011000001010000000011111001;
REG[2303] <= 32'b00000110000000100000011000000110;
REG[2304] <= 32'b11111001111111011111100100001101;
REG[2305] <= 32'b11111011111101101111001111100110;
REG[2306] <= 32'b00000000000011001111101011110001;
REG[2307] <= 32'b00000100000000111111110000001011;
REG[2308] <= 32'b00001011111111110000010011101110;
REG[2309] <= 32'b11110001000001100000111111111011;
REG[2310] <= 32'b00000010111110011110111100001101;
REG[2311] <= 32'b00001110111111111111110000001011;
REG[2312] <= 32'b00001100111011011111110011110111;
REG[2313] <= 32'b11101110000000011111111011101001;
REG[2314] <= 32'b11111001111011111110101011111111;
REG[2315] <= 32'b00000111110111101110110011101101;
REG[2316] <= 32'b11111101000001100001010111111001;
REG[2317] <= 32'b11110101000001001111001100000010;
REG[2318] <= 32'b00000101111110111111001111111011;
REG[2319] <= 32'b11110011111101011111110100000000;
REG[2320] <= 32'b00000011000001011111011111110011;
REG[2321] <= 32'b11111001000000111111101100000010;
REG[2322] <= 32'b11101100111011111111011011110001;
REG[2323] <= 32'b11101111111010111110100111110101;
REG[2324] <= 32'b11111010111101001110111011110110;
REG[2325] <= 32'b00000111000000100000111011111000;
REG[2326] <= 32'b00000111000011100000001111111011;
REG[2327] <= 32'b00000101111101101111010000000101;
REG[2328] <= 32'b11101110111011001111010100000010;
REG[2329] <= 32'b00000010111111111111101011110100;
REG[2330] <= 32'b11110111111100001111001011110111;
REG[2331] <= 32'b11101101111111101111111011110011;
REG[2332] <= 32'b11101110000000111110100011111010;
REG[2333] <= 32'b11111100000000011110101100001000;
REG[2334] <= 32'b11111001111111010001100011110100;
REG[2335] <= 32'b00000111111010100000111011111100;
REG[2336] <= 32'b11110010111110100001010100000001;
REG[2337] <= 32'b11111110111101001111101011110110;
REG[2338] <= 32'b00010010111111011111110111111100;
REG[2339] <= 32'b00000011111011111111000011110111;
REG[2340] <= 32'b11110000111101110000110011110000;
REG[2341] <= 32'b11101001111100100000001000010000;
REG[2342] <= 32'b00010001111100011101110111110011;
REG[2343] <= 32'b00000011111100111111001000001001;
REG[2344] <= 32'b11110111111100010000001111111011;
REG[2345] <= 32'b11110100000011011111100111101011;
REG[2346] <= 32'b00001100111111011111001000000100;
REG[2347] <= 32'b11111100111010001111101011101101;
REG[2348] <= 32'b11111000111101101111010111111111;
REG[2349] <= 32'b11111100111100111111011111110101;
REG[2350] <= 32'b11110110111111111111011011110111;
REG[2351] <= 32'b11111010111101101110101111110010;
REG[2352] <= 32'b11110011000000110000011011111000;
REG[2353] <= 32'b11110101111101101111111100001001;
REG[2354] <= 32'b00000111111110011111111011111010;
REG[2355] <= 32'b11111001000001100000010011111000;
REG[2356] <= 32'b00000011111111101111101011110110;
REG[2357] <= 32'b11111010111110011111110011110100;
REG[2358] <= 32'b11110110111101001111100100000011;
REG[2359] <= 32'b00000010111101101111011011110110;
REG[2360] <= 32'b11110111111111100000000111101011;
REG[2361] <= 32'b00000100111111110000001011111011;
REG[2362] <= 32'b11100010111010001111100100000100;
REG[2363] <= 32'b00101001110111101100110111010101;
REG[2364] <= 32'b00001000111111110000010100001110;
REG[2365] <= 32'b11111101000001111111111100000000;
REG[2366] <= 32'b00000101000000000000100000000111;
REG[2367] <= 32'b00000100111110110000000000001110;
REG[2368] <= 32'b00001111000101100000010000000011;
REG[2369] <= 32'b00000010000011101111010011101101;
REG[2370] <= 32'b11111100111101110000001100000110;
REG[2371] <= 32'b00001111000000111111101111111011;
REG[2372] <= 32'b00000011111100111110101011110011;
REG[2373] <= 32'b00001010111111010000100011111011;
REG[2374] <= 32'b11111001111011001111100000000010;
REG[2375] <= 32'b00000011111110111111011000000010;
REG[2376] <= 32'b00000011111110111111100111110111;
REG[2377] <= 32'b11110111000010000000100011111110;
REG[2378] <= 32'b11111001111110001111101000000000;
REG[2379] <= 32'b11110000111101101111111111111100;
REG[2380] <= 32'b11111011111110101111011011110111;
REG[2381] <= 32'b00000000111101001111100111111000;
REG[2382] <= 32'b11111101111110001111011111110101;
REG[2383] <= 32'b00000001111110011111111000000010;
REG[2384] <= 32'b00000101111110111111110100000001;
REG[2385] <= 32'b11111110111111110000001011111100;
REG[2386] <= 32'b00000101000011001111010000000000;
REG[2387] <= 32'b00001010111110111111100011111011;
REG[2388] <= 32'b00000101111110001111101011110100;
REG[2389] <= 32'b11111101000100010000100011101010;
REG[2390] <= 32'b11110010111110111110010111110100;
REG[2391] <= 32'b00000110111110101111011100001100;
REG[2392] <= 32'b00000111000010101110011111101010;
REG[2393] <= 32'b00000011000000001111110011111101;
REG[2394] <= 32'b11101100111011000000001011111110;
REG[2395] <= 32'b11110011111111100000001111111101;
REG[2396] <= 32'b00000100000001101111110000000001;
REG[2397] <= 32'b00001000000010000000110011111101;
REG[2398] <= 32'b00001001111100001111100011110010;
REG[2399] <= 32'b11110110000000000000001000001000;
REG[2400] <= 32'b11110101111101010000010011110010;
REG[2401] <= 32'b11110110111110101111111111111100;
REG[2402] <= 32'b11111110111111000000001011110110;
REG[2403] <= 32'b11111001111101101111101111101011;
REG[2404] <= 32'b11101111111100001111001011110011;
REG[2405] <= 32'b11110101000011000000011011110110;
REG[2406] <= 32'b11111011111111101111011100000101;
REG[2407] <= 32'b00000001000000101111101011110110;
REG[2408] <= 32'b11110111000011110000001100000011;
REG[2409] <= 32'b11110110111110011111010100000111;
REG[2410] <= 32'b00001111000011111111011011111100;
REG[2411] <= 32'b11111011000011110000001011111111;
REG[2412] <= 32'b11111011111111101111010100000011;
REG[2413] <= 32'b11111100111110111111110000000000;
REG[2414] <= 32'b11111000000001101111101111110100;
REG[2415] <= 32'b11111110111110101111110011111111;
REG[2416] <= 32'b11111111000001001111100100000100;
REG[2417] <= 32'b00000111111110111111101011111111;
REG[2418] <= 32'b11110011111110111111110100001000;
REG[2419] <= 32'b00000110111111100000110100010010;
REG[2420] <= 32'b11111111000010100000010011111000;
REG[2421] <= 32'b00010001000111100000110000001001;
REG[2422] <= 32'b00000011111101110000111000010010;
REG[2423] <= 32'b00000110000010000000010111111001;
REG[2424] <= 32'b00000000111101011111110000000100;
REG[2425] <= 32'b11111111000010010000100111110100;
REG[2426] <= 32'b11111100111101101111101111111011;
REG[2427] <= 32'b00000001111110100001010000000000;
REG[2428] <= 32'b00010001111110011111001111110100;
REG[2429] <= 32'b00000000111110011110111111111010;
REG[2430] <= 32'b11110101111100001111111000000001;
REG[2431] <= 32'b11101100111100011111011011111011;
REG[2432] <= 32'b11111111000011010000001011111010;
REG[2433] <= 32'b11110001000001010000111011111111;
REG[2434] <= 32'b00000011111110101111011100011010;
REG[2435] <= 32'b00011101000000000000001000000100;
REG[2436] <= 32'b11110011000010110001001100000001;
REG[2437] <= 32'b11111011000010011111001111111000;
REG[2438] <= 32'b11111011111111101111111100000000;
REG[2439] <= 32'b11101111111101101111011011111001;
REG[2440] <= 32'b11101110111110011111001011110100;
REG[2441] <= 32'b11111010000100010000001111111011;
REG[2442] <= 32'b11111001111101101111000000001000;
REG[2443] <= 32'b00001010111110111111111011110100;
REG[2444] <= 32'b11101001000010101111001011110010;
REG[2445] <= 32'b11110110111101101110111000001010;
REG[2446] <= 32'b00001111111101001110111111110010;
REG[2447] <= 32'b11110100111100011111101011111000;
REG[2448] <= 32'b11101110111100001111001111100111;
REG[2449] <= 32'b11100111111010001111101111111000;
REG[2450] <= 32'b11110111111010101110101011101010;
REG[2451] <= 32'b00001100000101100000110100001011;
REG[2452] <= 32'b00000000000000000000111100010101;
REG[2453] <= 32'b00001111111110011111011011110100;
REG[2454] <= 32'b00001010000001010000010100000101;
REG[2455] <= 32'b11111110111101111111101111111011;
REG[2456] <= 32'b11111111111011111111010011111010;
REG[2457] <= 32'b11111100000000000000001011111001;
REG[2458] <= 32'b11111001111101111111101111111101;
REG[2459] <= 32'b11111101111110001111110011111100;
REG[2460] <= 32'b11101001111110110000010111111001;
REG[2461] <= 32'b11111100000111011111000111110100;
REG[2462] <= 32'b00000001111111111110111100001010;
REG[2463] <= 32'b11101101000000010000100011111101;
REG[2464] <= 32'b11101000111100101111101111111110;
REG[2465] <= 32'b11111111111110101111110000000011;
REG[2466] <= 32'b11111100111101111111100111111001;
REG[2467] <= 32'b11111101000100011111100011110001;
REG[2468] <= 32'b11111000000001011111111100000011;
REG[2469] <= 32'b11110100111111101111110100011001;
REG[2470] <= 32'b00010100111101101111110111111110;
REG[2471] <= 32'b00001000111111110001000011111110;
REG[2472] <= 32'b11111110111111001111101111110111;
REG[2473] <= 32'b11110101111110100000101100000101;
REG[2474] <= 32'b00000101111111001111010111111011;
REG[2475] <= 32'b00000001111101111111101111110111;
REG[2476] <= 32'b11101011111100010000001011111010;
REG[2477] <= 32'b00000101111110111111001011111010;
REG[2478] <= 32'b11111111000011110000001000001110;
REG[2479] <= 32'b00000001111110111111000100001100;
REG[2480] <= 32'b00100000000001010000000111100011;
REG[2481] <= 32'b11110111000000010000111100010111;
REG[2482] <= 32'b00011000000001010000010111111101;
REG[2483] <= 32'b00000000111111000000001000000100;
REG[2484] <= 32'b11111010111111010000100100001100;
REG[2485] <= 32'b00010100000010100000000011111101;
REG[2486] <= 32'b00000101111111110001000000001010;
REG[2487] <= 32'b00001111111111000000010000001001;
REG[2488] <= 32'b00001010111111010000100011110101;
REG[2489] <= 32'b11111110000001110000000011110110;
REG[2490] <= 32'b00010110000000001111111100000010;
REG[2491] <= 32'b00000011111111000000000000000011;
REG[2492] <= 32'b11111111111111001111110100000101;
REG[2493] <= 32'b11111011111111111111110111111011;
REG[2494] <= 32'b11111000000001011111101100000000;
REG[2495] <= 32'b11111100111110001111100111111111;
REG[2496] <= 32'b00001011111101111111010111110111;
REG[2497] <= 32'b11111100111101110001101000000100;
REG[2498] <= 32'b11110101111111000000111011111110;
REG[2499] <= 32'b00010100000001011111001111110001;
REG[2500] <= 32'b11111101000000110000000111101110;
REG[2501] <= 32'b11110100111100001111111011110111;
REG[2502] <= 32'b00011110000000101111000011101101;
REG[2503] <= 32'b00000000111110110001011011110100;
REG[2504] <= 32'b11111101111110100000111011111011;
REG[2505] <= 32'b11111100000000111111110100001001;
REG[2506] <= 32'b11110111111010000001110000010101;
REG[2507] <= 32'b00010001000100101111010011101010;
REG[2508] <= 32'b00000100000000110000010111111000;
REG[2509] <= 32'b11110100000000100000000000010100;
REG[2510] <= 32'b00010011111111001111010100000010;
REG[2511] <= 32'b00000011111100011111101111111101;
REG[2512] <= 32'b11110001111111111111111100010000;
REG[2513] <= 32'b00010110000010010000000100001010;
REG[2514] <= 32'b11101110111101110000111100000000;
REG[2515] <= 32'b11110101111010010000001101001001;
REG[2516] <= 32'b11110110000001001110001111101111;
REG[2517] <= 32'b00000000001111100000110100010010;
REG[2518] <= 32'b11111100111100010000000011111101;
REG[2519] <= 32'b11111111111101111111011011110101;
REG[2520] <= 32'b11111011111011011111100100001010;
REG[2521] <= 32'b11111111000001101111110111111010;
REG[2522] <= 32'b11111110111100111111001111111011;
REG[2523] <= 32'b00000101000000110000011111111010;
REG[2524] <= 32'b11111101000001001111111111110100;
REG[2525] <= 32'b11111100111110101111100111111101;
REG[2526] <= 32'b11111001111110010000000100010010;
REG[2527] <= 32'b11111110000000000000001100001111;
REG[2528] <= 32'b00000100111010110000100000010110;
REG[2529] <= 32'b00100011000110011111111111110000;
REG[2530] <= 32'b11111110000111010000110000000011;
REG[2531] <= 32'b00000000111001101111010100010001;
REG[2532] <= 32'b00000101111010001111010000000111;
REG[2533] <= 32'b00110011111101111111110011101011;
REG[2534] <= 32'b11110111000101000001001011110011;
REG[2535] <= 32'b00000110111101110000101011110111;
REG[2536] <= 32'b11101010111100010000110000000010;
REG[2537] <= 32'b00001001111111001111100111110110;
REG[2538] <= 32'b00001100000001010000101000000000;
REG[2539] <= 32'b00000001111110010001100000001101;
REG[2540] <= 32'b00000110111100100001110000000001;
REG[2541] <= 32'b11110110111111000000001011111011;
REG[2542] <= 32'b00010111000100011110111011110101;
REG[2543] <= 32'b00000100111010100011100100100000;
REG[2544] <= 32'b11101011111011010000010011110111;
REG[2545] <= 32'b11110011111000011110111111111010;
REG[2546] <= 32'b11111000000011000000000011110001;
REG[2547] <= 32'b00100010111110111110111000100000;
REG[2548] <= 32'b00001010111100100001010111111001;
REG[2549] <= 32'b11110110111111111111111011111110;
REG[2550] <= 32'b00001100000100011110010011111100;
REG[2551] <= 32'b11101110111011100001101100011010;
REG[2552] <= 32'b11111101000001001110110011110000;
REG[2553] <= 32'b00001110000001111111101000010000;
REG[2554] <= 32'b11111110111111001111001011110001;
REG[2555] <= 32'b11110011111000100000100000000101;
REG[2556] <= 32'b00000100111111001111100011100001;
REG[2557] <= 32'b00010111000010101111001011111000;
REG[2558] <= 32'b11111001111101010000011011110101;
REG[2559] <= 32'b00000011111100010000011000000111;
REG[2560] <= 32'b00000011000001010000101100001001;
REG[2561] <= 32'b00000010000000111111111100010000;
REG[2562] <= 32'b00001000111111001111001100000011;
REG[2563] <= 32'b11111011111110000000110100000100;
REG[2564] <= 32'b00001101111110001111111100000000;
REG[2565] <= 32'b11111111111111001111111111111001;
REG[2566] <= 32'b00001000000010000000001100000110;
REG[2567] <= 32'b11111110111101101111111000000110;
REG[2568] <= 32'b11101111111111110000001100000110;
REG[2569] <= 32'b11111011000010011111101100100000;
REG[2570] <= 32'b00000111111110011111100000010100;
REG[2571] <= 32'b11111100000010011111010100000100;
REG[2572] <= 32'b11110110000000000000101000000010;
REG[2573] <= 32'b11111100111101010000000000001110;
REG[2574] <= 32'b00100101111111111111011111110100;
REG[2575] <= 32'b00001000001001000000000011110100;
REG[2576] <= 32'b00000101111010101111111100010111;
REG[2577] <= 32'b11111010111111111111010100010000;
REG[2578] <= 32'b11111111111000100000101100011110;
REG[2579] <= 32'b11110101000101101111101111011010;
REG[2580] <= 32'b00000010000001011111100100001100;
REG[2581] <= 32'b00000110000001010000001111111101;
REG[2582] <= 32'b00000010000010000000000011111001;
REG[2583] <= 32'b11111010111100111111010011110111;
REG[2584] <= 32'b11110111111101110000000100000010;
REG[2585] <= 32'b00000100000000000000001011111011;
REG[2586] <= 32'b00000000111111110000010011111101;
REG[2587] <= 32'b11111010111111010000010100000101;
REG[2588] <= 32'b00001000000000110001110100000010;
REG[2589] <= 32'b11110111111101010000001100000010;
REG[2590] <= 32'b00010011000100000000110011111110;
REG[2591] <= 32'b11111001111101011111100000000100;
REG[2592] <= 32'b00101000000010001111100100000111;
REG[2593] <= 32'b11111010111111000001000100000010;
REG[2594] <= 32'b11111011000000111111110011101001;
REG[2595] <= 32'b11110110111111010000010111111100;
REG[2596] <= 32'b00000100000000101111010000000011;
REG[2597] <= 32'b00001100111111101111001111111100;
REG[2598] <= 32'b00000100000000100000011100001000;
REG[2599] <= 32'b11111000000001001111100111111111;
REG[2600] <= 32'b00001101000010110000011000010011;
REG[2601] <= 32'b11110000111100111111011011111110;
REG[2602] <= 32'b11110010000000011111001011111011;
REG[2603] <= 32'b11111101111110111110110111101110;
REG[2604] <= 32'b00000011000100000001010000001111;
REG[2605] <= 32'b00001101111111111111111100010001;
REG[2606] <= 32'b00000010000010110000010100000010;
REG[2607] <= 32'b00000110000010010000011100000100;
REG[2608] <= 32'b00100000111011011111001000000001;
REG[2609] <= 32'b00000100111111011111001011110110;
REG[2610] <= 32'b11101001111100111111100011111010;
REG[2611] <= 32'b11101101111110011110101111110111;
REG[2612] <= 32'b11111101000011011111101011111001;
REG[2613] <= 32'b11110000111101011110111011111110;
REG[2614] <= 32'b11110111000001100000100111111110;
REG[2615] <= 32'b11110111111110001111101111111101;
REG[2616] <= 32'b00010011111111101111000000000001;
REG[2617] <= 32'b11111100000101001111101011111101;
REG[2618] <= 32'b00001001111111011111101100010010;
REG[2619] <= 32'b00000110111111000000010111110110;
REG[2620] <= 32'b11110011000011010000010111111111;
REG[2621] <= 32'b00001001111101011110111100001000;
REG[2622] <= 32'b11111100111110111110011000001000;
REG[2623] <= 32'b00010000000110001110111011101100;
REG[2624] <= 32'b11100101000101110000111100010010;
REG[2625] <= 32'b11101100111101101110110000000001;
REG[2626] <= 32'b00000000000000101111110111111111;
REG[2627] <= 32'b11110111000000011111000111101100;
REG[2628] <= 32'b00001000111101001111000000010000;
REG[2629] <= 32'b11111110111101001111111011111111;
REG[2630] <= 32'b11110101111011111110111011101011;
REG[2631] <= 32'b00000110000000000000100111110110;
REG[2632] <= 32'b00000110000001111110111011110111;
REG[2633] <= 32'b00000101000001110001000000010000;
REG[2634] <= 32'b11111010000011010001100011111010;
REG[2635] <= 32'b11111011111110110001000000000001;
REG[2636] <= 32'b00000001111101101111100100000110;
REG[2637] <= 32'b00011010000101001111101111110111;
REG[2638] <= 32'b11110111111111010001010100001111;
REG[2639] <= 32'b00000011111011001111011100000101;
REG[2640] <= 32'b11110110111111111111111000001100;
REG[2641] <= 32'b11111101000000011111011011111111;
REG[2642] <= 32'b00001110000101000000100100001010;
REG[2643] <= 32'b11110001111111011111111100011000;
REG[2644] <= 32'b00000010111101111111111000000100;
REG[2645] <= 32'b00000011111110110000001111111101;
REG[2646] <= 32'b11110111000001111111101000001001;
REG[2647] <= 32'b00001111000000001111011000001000;
REG[2648] <= 32'b00000011000001000000010011111100;
REG[2649] <= 32'b11110101000011010000111111111100;
REG[2650] <= 32'b11111111111111001111111100000101;
REG[2651] <= 32'b00001001000101001111011000001011;
REG[2652] <= 32'b11111110000110010000010111111111;
REG[2653] <= 32'b11110110000001111111110000000100;
REG[2654] <= 32'b00001011111010111111100000000010;
REG[2655] <= 32'b11110111111110110000101111101010;
REG[2656] <= 32'b11101001111100101111010000000001;
REG[2657] <= 32'b00000100111110101111010000000001;
REG[2658] <= 32'b00000011000010111111110111111010;
REG[2659] <= 32'b00000010000000101111110100000011;
REG[2660] <= 32'b11110110111110101111101000000110;
REG[2661] <= 32'b11111011000010001111101111111011;
REG[2662] <= 32'b11110101000011101111001111111001;
REG[2663] <= 32'b11111110000101010001001100001000;
REG[2664] <= 32'b11110011000000111111111000011000;
REG[2665] <= 32'b00010010000001011110101100000000;
REG[2666] <= 32'b11111110000100100001001000000001;
REG[2667] <= 32'b11111001111101111111101000001010;
REG[2668] <= 32'b11110111000101111111101000000000;
REG[2669] <= 32'b11110111000000000000001000001111;
REG[2670] <= 32'b11110100111111001111110011111001;
REG[2671] <= 32'b00000011000010001111011000001110;
REG[2672] <= 32'b00000111000100110001010000001101;
REG[2673] <= 32'b00000001000010110000010000000011;
REG[2674] <= 32'b00001001000011001111101100001101;
REG[2675] <= 32'b11111100111111111111111000000111;
REG[2676] <= 32'b00010000000001000000010100001001;
REG[2677] <= 32'b00000110000001011111010111111101;
REG[2678] <= 32'b00000001000101110000111111111011;
REG[2679] <= 32'b00001011000000110000011000001010;
REG[2680] <= 32'b11111111000000111111011000001100;
REG[2681] <= 32'b00001000000011110000000011101111;
REG[2682] <= 32'b11111011001010110001001000001110;
REG[2683] <= 32'b00000010111110101111110011111000;
REG[2684] <= 32'b00000001111100011111001011111111;
REG[2685] <= 32'b00001110000000010000010111111111;
REG[2686] <= 32'b00000011111111101111000011110101;
REG[2687] <= 32'b11110100111111101111001111101111;
REG[2688] <= 32'b11110110111100111111101011110111;
REG[2689] <= 32'b11101101111101001111011000000000;
REG[2690] <= 32'b00000001000011111111011111110101;
REG[2691] <= 32'b00000011000001100000010100000101;
REG[2692] <= 32'b00001010111100011110110011111000;
REG[2693] <= 32'b00000001111110011111010011110101;
REG[2694] <= 32'b00010010111100101111000111110100;
REG[2695] <= 32'b11111101111101000000100011101100;
REG[2696] <= 32'b11110000111111110000110000000010;
REG[2697] <= 32'b00001110111110001111101111110011;
REG[2698] <= 32'b00000101111111111111000111111101;
REG[2699] <= 32'b00001000000001000000100100000011;
REG[2700] <= 32'b11111001000000000000010011110110;
REG[2701] <= 32'b00000100000001001110011111110110;
REG[2702] <= 32'b11111110111101111111011011111001;
REG[2703] <= 32'b00000110000010000001000011101111;
REG[2704] <= 32'b11101101111100000000010100001110;
REG[2705] <= 32'b00011011111100111110110111110011;
REG[2706] <= 32'b00000100000011110001100011110111;
REG[2707] <= 32'b11110000111100011110110111110001;
REG[2708] <= 32'b11111101000010110000010011111011;
REG[2709] <= 32'b11101000111011111111101100001110;
REG[2710] <= 32'b00010100111111001111001011110100;
REG[2711] <= 32'b11111100000001000000101000001001;
REG[2712] <= 32'b00000001111110000000101011111001;
REG[2713] <= 32'b11101100000001111111010111110100;
REG[2714] <= 32'b11111111111110001110001111101001;
REG[2715] <= 32'b11111110111111100000010111110101;
REG[2716] <= 32'b11100110111110111111100000000010;
REG[2717] <= 32'b00001010000100000000100011111010;
REG[2718] <= 32'b00000010000110101111101100010001;
REG[2719] <= 32'b00000011111101110000001100000010;
REG[2720] <= 32'b11111101000001111111111100000000;
REG[2721] <= 32'b11111011111110001111100100001110;
REG[2722] <= 32'b00000001111111111111100111111101;
REG[2723] <= 32'b11111001111111111111101100000001;
REG[2724] <= 32'b11111011111111011111110011111110;
REG[2725] <= 32'b00000000111110111111101111110011;
REG[2726] <= 32'b11111100000011000000000011111010;
REG[2727] <= 32'b11110101111110011111110000000001;
REG[2728] <= 32'b11110011111101101111101100000000;
REG[2729] <= 32'b00000010111100001111100011111001;
REG[2730] <= 32'b11110011000000111111101111111001;
REG[2731] <= 32'b11101100111100001111011000000001;
REG[2732] <= 32'b11110001000000111111100111111001;
REG[2733] <= 32'b00000101000000011111010000000000;
REG[2734] <= 32'b11111111000000001110110111110000;
REG[2735] <= 32'b11111011000010001111111100000110;
REG[2736] <= 32'b11110110111111011111010000011000;
REG[2737] <= 32'b00000000000000011111110111111111;
REG[2738] <= 32'b11110100111111111111101111110111;
REG[2739] <= 32'b00000010000010000000001111110110;
REG[2740] <= 32'b11111010111101100000000000001011;
REG[2741] <= 32'b00001000111011001111011011111010;
REG[2742] <= 32'b00001110000100010001010111101010;
REG[2743] <= 32'b11101101111101000000001111111011;
REG[2744] <= 32'b00000011000011001111100100000010;
REG[2745] <= 32'b00001001111101000000100100001001;
REG[2746] <= 32'b00000111111110100000011111111011;
REG[2747] <= 32'b00001000000001100000000000000101;
REG[2748] <= 32'b00000000111110101111100111111010;
REG[2749] <= 32'b11110101000000001111100011011011;
REG[2750] <= 32'b11101101111100111111101000000011;
REG[2751] <= 32'b00000010111110011111111011110010;
REG[2752] <= 32'b11110110111110010000110111111011;
REG[2753] <= 32'b11111010000001010000111000000011;
REG[2754] <= 32'b00100111000010001111101000001001;
REG[2755] <= 32'b00001011000001111111100100001011;
REG[2756] <= 32'b00000010111111111111100100000101;
REG[2757] <= 32'b11111010111111010000000011101011;
REG[2758] <= 32'b11111101000000111111111011111100;
REG[2759] <= 32'b11110111111111001111110111111001;
REG[2760] <= 32'b11110010111100111111010111110101;
REG[2761] <= 32'b11111111000001001111100000000100;
REG[2762] <= 32'b00011010000001101111011000000011;
REG[2763] <= 32'b11110110111110100000111000000010;
REG[2764] <= 32'b00001001000011001111100000000001;
REG[2765] <= 32'b00000100111111110000000100011110;
REG[2766] <= 32'b00000110000000001111100111111011;
REG[2767] <= 32'b00001001111110101111101111111010;
REG[2768] <= 32'b11111000111110100000010111111100;
REG[2769] <= 32'b11111010111101011111101100000111;
REG[2770] <= 32'b00001011000001101111000000000100;
REG[2771] <= 32'b00000111000000000000101111111111;
REG[2772] <= 32'b11101100111101101111100011111000;
REG[2773] <= 32'b00001001000000011111011111110111;
REG[2774] <= 32'b11101110000000010000010000000001;
REG[2775] <= 32'b00000100111110001111011100001011;
REG[2776] <= 32'b11111111111110101111110111111000;
REG[2777] <= 32'b11111000111101101111111111111000;
REG[2778] <= 32'b00000010111111111111101100001010;
REG[2779] <= 32'b11111011111110111111011011110101;
REG[2780] <= 32'b11110100111111101111111011111011;
REG[2781] <= 32'b11110000111010111111000000001000;
REG[2782] <= 32'b00000010111100110000010111110111;
REG[2783] <= 32'b11111000111111111111011111110110;
REG[2784] <= 32'b00001100000011110000010011111110;
REG[2785] <= 32'b11110101111101111111110100001011;
REG[2786] <= 32'b11111011111100111111010111111101;
REG[2787] <= 32'b11111111000010011111110011110101;
REG[2788] <= 32'b11111100111100110000101011111100;
REG[2789] <= 32'b11111001000001100000010111110101;
REG[2790] <= 32'b00001011111111011111000100000000;
REG[2791] <= 32'b11111000111100010000010011111011;
REG[2792] <= 32'b11111010000000001111100111110110;
REG[2793] <= 32'b11111100111101101111110111111001;
REG[2794] <= 32'b11111101111110100000000111110011;
REG[2795] <= 32'b11110001111101100010101100111000;
REG[2796] <= 32'b00000011111101011111010011101111;
REG[2797] <= 32'b00000111000010011110101111101110;
REG[2798] <= 32'b11110000111100111111010111111110;
REG[2799] <= 32'b00001110111110011111010011111001;
REG[2800] <= 32'b11110011000000111111100011110010;
REG[2801] <= 32'b11110101111101111111011111111101;
REG[2802] <= 32'b00010100000001110000010111111011;
REG[2803] <= 32'b00000010000001000000100111111010;
REG[2804] <= 32'b00000001111110011111111111111011;
REG[2805] <= 32'b00000101111111110000000111110111;
REG[2806] <= 32'b11110111111101000000010011111111;
REG[2807] <= 32'b00000101000010000000000100000001;
REG[2808] <= 32'b11111101111110011111001111110111;
REG[2809] <= 32'b11101100111101100000000111111100;
REG[2810] <= 32'b11110111000011011111110011111100;
REG[2811] <= 32'b11110101111110001111100011111110;
REG[2812] <= 32'b11110011111110010000011000000011;
REG[2813] <= 32'b11111001111110001111011111111111;
REG[2814] <= 32'b11110111111111001111100111111011;
REG[2815] <= 32'b11111001111101111111000111111100;
REG[2816] <= 32'b00000110000001000000100100010101;
REG[2817] <= 32'b11111101000001001111111000000100;
REG[2818] <= 32'b00001010000100010000110000001100;
REG[2819] <= 32'b00000111111111110000000011111111;
REG[2820] <= 32'b00001000000000111110111011111101;
REG[2821] <= 32'b11111000000010000000011011111000;
REG[2822] <= 32'b11110100111100111111100000010001;
REG[2823] <= 32'b00000111000000110000011011111101;
REG[2824] <= 32'b00000001000010101110111100000010;
REG[2825] <= 32'b00000110000001011111010011111011;
REG[2826] <= 32'b11011110111011010000011011111110;
REG[2827] <= 32'b11101011111101011111100011111111;
REG[2828] <= 32'b00001100000001011111100100000101;
REG[2829] <= 32'b11111000111110111111101111110010;
REG[2830] <= 32'b11111100111110111111010111110000;
REG[2831] <= 32'b11110100111101101111011011111001;
REG[2832] <= 32'b00001100111110001111111011111101;
REG[2833] <= 32'b00000000000000000000100100001110;
REG[2834] <= 32'b11111110000000101111111000001000;
REG[2835] <= 32'b00000110111110000000110000000101;
REG[2836] <= 32'b11111011111110011111010011111111;
REG[2837] <= 32'b00000110000010011111100011111001;
REG[2838] <= 32'b11111010111100011111100000000110;
REG[2839] <= 32'b11111101000010101111100011101101;
REG[2840] <= 32'b11110110000000001111000000001010;
REG[2841] <= 32'b11111101111100011111111111111000;
REG[2842] <= 32'b11111010000011101111110011111010;
REG[2843] <= 32'b11110011111110110000011011110010;
REG[2844] <= 32'b00000011000001000000000111111001;
REG[2845] <= 32'b00000111111101110000001100000110;
REG[2846] <= 32'b11111010111110010000001111111010;
REG[2847] <= 32'b11111011111101101111010000010010;
REG[2848] <= 32'b00010010000010011111100111101111;
REG[2849] <= 32'b11111000000010110000011100000101;
REG[2850] <= 32'b11111100111110011111110100000111;
REG[2851] <= 32'b00001100000101001110111111110101;
REG[2852] <= 32'b11110001000010000000100100000001;
REG[2853] <= 32'b11111100000010101111011111111001;
REG[2854] <= 32'b00000101000001001111101100001001;
REG[2855] <= 32'b11111010111110000000001000000110;
REG[2856] <= 32'b00000000111101101111111100001000;
REG[2857] <= 32'b11110110111110101111110111110110;
REG[2858] <= 32'b11110101000001101111010011111011;
REG[2859] <= 32'b00001010000010010000010000001111;
REG[2860] <= 32'b11110011111111010001001100010010;
REG[2861] <= 32'b00001000111101111111111011111101;
REG[2862] <= 32'b00000011000101110000011011110100;
REG[2863] <= 32'b11110110111110111111000111111101;
REG[2864] <= 32'b00001001111100101111001011110111;
REG[2865] <= 32'b00000011111111111111011111111010;
REG[2866] <= 32'b11111001000001111111011100000010;
REG[2867] <= 32'b11111010000001100000010100001110;
REG[2868] <= 32'b00000000000100101111111111111001;
REG[2869] <= 32'b00000101000011100001000000000101;
REG[2870] <= 32'b00000011111110111111000111110111;
REG[2871] <= 32'b11111010111110001111100011110111;
REG[2872] <= 32'b11101101111110001111101111111010;
REG[2873] <= 32'b11111011000000101111101011111001;
REG[2874] <= 32'b01001001111111011111000011111111;
REG[2875] <= 32'b11111100111101000011001100001100;
REG[2876] <= 32'b11111010111101011111001111111000;
REG[2877] <= 32'b00000001000001011111101111110101;
REG[2878] <= 32'b11110100111110100000000111110010;
REG[2879] <= 32'b11111001111110001111011111110110;
REG[2880] <= 32'b00001000000000000000011111110011;
REG[2881] <= 32'b11110101111110010000011000001100;
REG[2882] <= 32'b00000001111111111111101111111010;
REG[2883] <= 32'b11111101000000110000110011110010;
REG[2884] <= 32'b11110101111101000000101000001010;
REG[2885] <= 32'b00001010000010110000100100001011;
REG[2886] <= 32'b00000110000011011111111000000011;
REG[2887] <= 32'b11111110000000011111010000000001;
REG[2888] <= 32'b00000000000011000001010100001000;
REG[2889] <= 32'b11111001111110101111101100000110;
REG[2890] <= 32'b00001000111111011111100111111100;
REG[2891] <= 32'b00000000111011010000001111111111;
REG[2892] <= 32'b00000110000000000000011011111100;
REG[2893] <= 32'b11111100000001010000001111111011;
REG[2894] <= 32'b00000000111110101111110111111111;
REG[2895] <= 32'b00000101111111111111101111111110;
REG[2896] <= 32'b00000011111110100000001011111111;
REG[2897] <= 32'b00001011111111110000111100001100;
REG[2898] <= 32'b11111101111110000000010100000000;
REG[2899] <= 32'b00001101000011101111111011111100;
REG[2900] <= 32'b00001011111111100000010100001100;
REG[2901] <= 32'b11110001000000101111110011110110;
REG[2902] <= 32'b11111011000001101111100011110001;
REG[2903] <= 32'b11111111000000100000010000001101;
REG[2904] <= 32'b11111101000000010000101100000111;
REG[2905] <= 32'b00000111000111101111111011110001;
REG[2906] <= 32'b11110110111111010000001100001011;
REG[2907] <= 32'b11111000111100110000001011110010;
REG[2908] <= 32'b00000010000100111111000011110001;
REG[2909] <= 32'b11111111111101110000000000001101;
REG[2910] <= 32'b00000100111111000000001000000000;
REG[2911] <= 32'b00000010111101110000000111110110;
REG[2912] <= 32'b11111110111111010001000000010111;
REG[2913] <= 32'b11111101111110100000100011110100;
REG[2914] <= 32'b00001011000101010000101011111011;
REG[2915] <= 32'b11110110000000000000001011110011;
REG[2916] <= 32'b11111100111110000000011111111110;
REG[2917] <= 32'b00000100111100111111111111110111;
REG[2918] <= 32'b00001000111101011111101111101111;
REG[2919] <= 32'b00011111000010010000010000000110;
REG[2920] <= 32'b11111110111111110000010111111001;
REG[2921] <= 32'b11111101000000111111010111111001;
REG[2922] <= 32'b00000011111101011111111000000110;
REG[2923] <= 32'b11111100000000010000111100001100;
REG[2924] <= 32'b00000000111111110000011100010100;
REG[2925] <= 32'b00010001000010010000011111111011;
REG[2926] <= 32'b00000100000101010001001000001011;
REG[2927] <= 32'b00000110111110010000001000001010;
REG[2928] <= 32'b00010110111110111110110011111000;
REG[2929] <= 32'b11110111111100010000111000001001;
REG[2930] <= 32'b11111010111110011111110011110110;
REG[2931] <= 32'b00001000000010001111000000000100;
REG[2932] <= 32'b00010111000010100001000000010011;
REG[2933] <= 32'b00000101111111100000100100000111;
REG[2934] <= 32'b01000000000111101111110111110010;
REG[2935] <= 32'b00000101000001100000100100001011;
REG[2936] <= 32'b00000011000010010000001100001011;
REG[2937] <= 32'b11111100111111100000000011111001;
REG[2938] <= 32'b11110111111111000000010100001110;
REG[2939] <= 32'b00000100111010001110100011111011;
REG[2940] <= 32'b00001000000001110000010111101110;
REG[2941] <= 32'b11111001000010100000110000000000;
REG[2942] <= 32'b00010111000010100001001000001001;
REG[2943] <= 32'b00011010000001000011001000001010;
REG[2944] <= 32'b00011100000000110000000000000101;
REG[2945] <= 32'b00000101111111100000101000000100;
REG[2946] <= 32'b00000111111110011111011011110100;
REG[2947] <= 32'b11111010000000100001001000000110;
REG[2948] <= 32'b00000000111101011111100100100010;
REG[2949] <= 32'b00001001000010000000011111101110;
REG[2950] <= 32'b00100001001111001111001011110111;
REG[2951] <= 32'b00001010000010110001000111110111;
REG[2952] <= 32'b11101010111100110000000100110010;
REG[2953] <= 32'b00101010000000101110100111110010;
REG[2954] <= 32'b00000000000011100001111011111111;
REG[2955] <= 32'b11111010111110011111011000000111;
REG[2956] <= 32'b00001011000011001111101011111110;
REG[2957] <= 32'b11101110111111110000000000000000;
REG[2958] <= 32'b11110101111100101110101011110101;
REG[2959] <= 32'b00000000000001000000010000000110;
REG[2960] <= 32'b00001010000000111111010111111001;
REG[2961] <= 32'b00000010000001010000011000000010;
REG[2962] <= 32'b11110001111101011111110100000111;
REG[2963] <= 32'b00001001000011111111110111111011;
REG[2964] <= 32'b11101111111010111111100011110011;
REG[2965] <= 32'b11101100111101001111010011111011;
REG[2966] <= 32'b11111111111110011111001100001001;
REG[2967] <= 32'b11110000111100101111101011111100;
REG[2968] <= 32'b00000001000101000010110000011110;
REG[2969] <= 32'b11101011000000010001100111111101;
REG[2970] <= 32'b00111011001001001110001100001010;
REG[2971] <= 32'b00100010111111011110110011111000;
REG[2972] <= 32'b11011111000010010000011011111111;
REG[2973] <= 32'b00000001111110000000001100000110;
REG[2974] <= 32'b11110110111111101111000111101011;
REG[2975] <= 32'b11110001000010110000000100000001;
REG[2976] <= 32'b11101100111100001111100011110111;
REG[2977] <= 32'b11111100000001011111010100000001;
REG[2978] <= 32'b00000101111111010000110100000000;
REG[2979] <= 32'b11111110000111000001000000011000;
REG[2980] <= 32'b00010111000000111111001000001011;
REG[2981] <= 32'b00000000000000100000101100000101;
REG[2982] <= 32'b11111100111111001111001100000000;
REG[2983] <= 32'b00001011000010101111100111111000;
REG[2984] <= 32'b11110010111111100000001000001000;
REG[2985] <= 32'b11111011111101011111100000001000;
REG[2986] <= 32'b11111101000001001111010011110111;
REG[2987] <= 32'b11110101000100000000010100001011;
REG[2988] <= 32'b11110010111100111111010100001100;
REG[2989] <= 32'b00000111111111101111101011110101;
REG[2990] <= 32'b11110011000010010000011000001011;
REG[2991] <= 32'b00000110111111110000001111110001;
REG[2992] <= 32'b11110110111101001111111111110010;
REG[2993] <= 32'b11111011111100001111100111110011;
REG[2994] <= 32'b00000010000000000000100011100111;
REG[2995] <= 32'b00000000111110001111101111110000;
REG[2996] <= 32'b11101100000100100000100000001001;
REG[2997] <= 32'b11110011111101011111000000001111;
REG[2998] <= 32'b00000000000010011111011011111001;
REG[2999] <= 32'b11110101000010010000100000001010;
REG[3000] <= 32'b11110011111101111111111111111011;
REG[3001] <= 32'b00001010000100000000010000000111;
REG[3002] <= 32'b11111011111011111111101000001001;
REG[3003] <= 32'b11111000111011101110111000001010;
REG[3004] <= 32'b11110111111011010000011100000110;
REG[3005] <= 32'b11110101000001010001111100001000;
REG[3006] <= 32'b11111110000000101110110100001110;
REG[3007] <= 32'b00101101000011000000010000000011;
REG[3008] <= 32'b11110010111110010001100111110011;
REG[3009] <= 32'b00011101001000000000101100000101;
REG[3010] <= 32'b00000000000001011111100100000000;
REG[3011] <= 32'b11111100000000011111010100000101;
REG[3012] <= 32'b11111011000000101111011000001001;
REG[3013] <= 32'b00000011000001100000001111111101;
REG[3014] <= 32'b00000000000000000001111000000001;
REG[3015] <= 32'b11111101111111111111100100011011;
REG[3016] <= 32'b00110010000100110000000011111010;
REG[3017] <= 32'b11111110000001000011010000001000;
REG[3018] <= 32'b11011101111000101110110100000010;
REG[3019] <= 32'b00000111000101001110011011101001;
REG[3020] <= 32'b11100111111111000000000100010001;
REG[3021] <= 32'b11111001111110011111010000000100;
REG[3022] <= 32'b00001001000000111111100111111110;
REG[3023] <= 32'b00001110000001000001001100010011;
REG[3024] <= 32'b11110111111111100000111000011001;
REG[3025] <= 32'b00010000000011001111110100000001;
REG[3026] <= 32'b00000010000010100000010000000000;
REG[3027] <= 32'b00001101000011010000111011110001;
REG[3028] <= 32'b11110001000000000001100100001110;
REG[3029] <= 32'b00001100000011101111110111111110;
REG[3030] <= 32'b00010000000010100000010100001010;
REG[3031] <= 32'b11111111111111101110111011111001;
REG[3032] <= 32'b00000011000101111111110011101110;
REG[3033] <= 32'b11101110111101100000000100110010;
REG[3034] <= 32'b00000100111100101111000011110010;
REG[3035] <= 32'b11111000000110110000010111111100;
REG[3036] <= 32'b00000100111110011111100111110011;
REG[3037] <= 32'b11111001111101110000010100001100;
REG[3038] <= 32'b00000100111101111111111111110100;
REG[3039] <= 32'b11111110111111101111101011110000;
REG[3040] <= 32'b11110111111101011111001111101110;
REG[3041] <= 32'b11110010000100001111111000010110;
REG[3042] <= 32'b11111100111101111111010000010110;
REG[3043] <= 32'b00000001000000001111101011111001;
REG[3044] <= 32'b11111101000101010001011000010111;
REG[3045] <= 32'b11111111111111010000000100000101;
REG[3046] <= 32'b00001111000001111111010111110110;
REG[3047] <= 32'b00000010000001100000011100000011;
REG[3048] <= 32'b11101111111111010000101111110010;
REG[3049] <= 32'b00000101111111011111110011110000;
REG[3050] <= 32'b11110100000011110000011100001000;
REG[3051] <= 32'b00000001111101111111110000000111;
REG[3052] <= 32'b11111101111110011111011111111011;
REG[3053] <= 32'b00000110000000110000001011111001;
REG[3054] <= 32'b00010010000010100000100000000110;
REG[3055] <= 32'b11111111000000010001111011110110;
REG[3056] <= 32'b11111000111111001111001011110100;
REG[3057] <= 32'b00011001111110011111110011110000;
REG[3058] <= 32'b11110000111100111111110111111101;
REG[3059] <= 32'b00000111000001100000101100001110;
REG[3060] <= 32'b11111000111101110000010000011100;
REG[3061] <= 32'b00111111000100101111110000000100;
REG[3062] <= 32'b11111110000001000001010100000100;
REG[3063] <= 32'b00001100000110100001000100001000;
REG[3064] <= 32'b11111111000011010000010100010001;
REG[3065] <= 32'b00000001111111001111011111110011;
REG[3066] <= 32'b11111001000010001111100011111001;
REG[3067] <= 32'b11110011111111001110011111110110;
REG[3068] <= 32'b11111110000011100010000000010100;
REG[3069] <= 32'b11101000111101000000101100000010;
REG[3070] <= 32'b00001111000101001110111111101000;
REG[3071] <= 32'b00001110000001000000110000001001;
REG[3072] <= 32'b11111110000001100000010100101010;
REG[3073] <= 32'b00000101000000010000000000001010;
REG[3074] <= 32'b00000101000100010000000100000100;
REG[3075] <= 32'b11111101111110110000000000001011;
REG[3076] <= 32'b11110111000011110000010100001001;
REG[3077] <= 32'b00000000000010111111001111111010;
REG[3078] <= 32'b00000110111111101111101000000011;
REG[3079] <= 32'b11110111000001001111111111111011;
REG[3080] <= 32'b00000010111111000000010100001100;
REG[3081] <= 32'b00000101111111111111110100001011;
REG[3082] <= 32'b00000100000001100001010000000101;
REG[3083] <= 32'b00000011000001111111110000000100;
REG[3084] <= 32'b11111101000000100000001111111101;
REG[3085] <= 32'b00001101000010000000010111110010;
REG[3086] <= 32'b11111110111110101111010100001110;
REG[3087] <= 32'b00001010111110000000101011110111;
REG[3088] <= 32'b00000001111110001111110011111100;
REG[3089] <= 32'b11111101000110100010000000000110;
REG[3090] <= 32'b11111101000000110000111100000110;
REG[3091] <= 32'b00000000111111101111001111110101;
REG[3092] <= 32'b00000001111111111111100000000110;
REG[3093] <= 32'b00001001000001000000011100000011;
REG[3094] <= 32'b00000000111101110000100111111111;
REG[3095] <= 32'b11111110000011110000100100000001;
REG[3096] <= 32'b00000000111101001111101100000000;
REG[3097] <= 32'b11111000111100110000001011111011;
REG[3098] <= 32'b11111111111110011110110011110011;
REG[3099] <= 32'b11110011111110101111111100000111;
REG[3100] <= 32'b11111101000000011110101111110011;
REG[3101] <= 32'b11110111000000110000010111110001;
REG[3102] <= 32'b11110111111101011111001100001000;
REG[3103] <= 32'b11111101111100100000110100010011;
REG[3104] <= 32'b00000111000010001111110011111011;
REG[3105] <= 32'b00011101000010010000010100000000;
REG[3106] <= 32'b11111110000010010000100011111101;
REG[3107] <= 32'b11111100111100111110111111110011;
REG[3108] <= 32'b00000010000000110000001000000110;
REG[3109] <= 32'b11110110000000011111101000000001;
REG[3110] <= 32'b11110111111111101111111000001010;
REG[3111] <= 32'b11110101111100111111100000001000;
REG[3112] <= 32'b00000101000000101111001011110111;
REG[3113] <= 32'b00001110000100001111111100000100;
REG[3114] <= 32'b11110110111111100001010111111000;
REG[3115] <= 32'b11110101000000010000110100001110;
REG[3116] <= 32'b00001111000000010000100000001000;
REG[3117] <= 32'b00000101000001110000000011111111;
REG[3118] <= 32'b11111001111110010000010000100011;
REG[3119] <= 32'b00101001000001111111001111110101;
REG[3120] <= 32'b11111000111110010000011000010100;
REG[3121] <= 32'b11111110111111011110011111101111;
REG[3122] <= 32'b00000011000111101111110111110000;
REG[3123] <= 32'b11100110111010110000001000001110;
REG[3124] <= 32'b11111100111111011110110111111001;
REG[3125] <= 32'b00001011111011011110101011111110;
REG[3126] <= 32'b11110111111110011111011100000001;
REG[3127] <= 32'b00000010000000101111001111111110;
REG[3128] <= 32'b11111000111111100000001111111100;
REG[3129] <= 32'b11111000111111001111010011110111;
REG[3130] <= 32'b11111010111110001111101111101011;
REG[3131] <= 32'b11110100111110101111111100000000;
REG[3132] <= 32'b11110111111011011111011111111010;
REG[3133] <= 32'b00000000000010110000001000000000;
REG[3134] <= 32'b00000000111110011111110000001100;
REG[3135] <= 32'b00000011000011100000010100000001;
REG[3136] <= 32'b11111101111100000000000000000001;
REG[3137] <= 32'b11111100000001100000011000000100;
REG[3138] <= 32'b00000101000000011111100100000100;
REG[3139] <= 32'b00000101000001010000001100010100;
REG[3140] <= 32'b00000100111001111111010011111011;
REG[3141] <= 32'b00001100000100110000001011111100;
REG[3142] <= 32'b11110101000010000000101100001001;
REG[3143] <= 32'b00000111111101100000010000001101;
REG[3144] <= 32'b00000000000010000000011011110011;
REG[3145] <= 32'b11110111111111010000011100001101;
REG[3146] <= 32'b00011001111110111111001011111101;
REG[3147] <= 32'b11111100000001000000001000000011;
REG[3148] <= 32'b11110001000000101110111111110111;
REG[3149] <= 32'b11111010000110001111000011100100;
REG[3150] <= 32'b11110011111111110000011100000001;
REG[3151] <= 32'b11110001111110000000011100000011;
REG[3152] <= 32'b00000110111011101110111000000011;
REG[3153] <= 32'b00010101000010010000000000001000;
REG[3154] <= 32'b11110111111100110001011000010101;
REG[3155] <= 32'b00000011000001101111100111110010;
REG[3156] <= 32'b00000100000010011111011100000100;
REG[3157] <= 32'b11111101000010101111111100000011;
REG[3158] <= 32'b00001010000011111111100111110010;
REG[3159] <= 32'b11101010111101010000010011111111;
REG[3160] <= 32'b11110111111110001111010011111101;
REG[3161] <= 32'b00001101111010111111011111110101;
REG[3162] <= 32'b11111010111111001111100111111100;
REG[3163] <= 32'b00000111000000100000010100001110;
REG[3164] <= 32'b00001000111110100000010000001100;
REG[3165] <= 32'b11111100000000101111100100000100;
REG[3166] <= 32'b00000001000000111111100000001010;
REG[3167] <= 32'b11111100000001110000100111110100;
REG[3168] <= 32'b00001111000100111111100100000110;
REG[3169] <= 32'b11110101111101000000010100000101;
REG[3170] <= 32'b11111100111100011110100111111001;
REG[3171] <= 32'b00001111000000100000001000000111;
REG[3172] <= 32'b00001100000000100000000011111101;
REG[3173] <= 32'b11111101111110110000000011111010;
REG[3174] <= 32'b00001100000010000001011100000110;
REG[3175] <= 32'b00000010111101101111101011110111;
REG[3176] <= 32'b11111011111101100000001111111111;
REG[3177] <= 32'b11111110111110101111111011111011;
REG[3178] <= 32'b00000100000010001111010111110001;
REG[3179] <= 32'b11111001111111111111100100000110;
REG[3180] <= 32'b00000011111010101111001111111011;
REG[3181] <= 32'b00001010000001110000011000000010;
REG[3182] <= 32'b00000011000001000000100000001010;
REG[3183] <= 32'b00001000111110100000100011111101;
REG[3184] <= 32'b11111101000001000000000000000010;
REG[3185] <= 32'b00001000111110101111111111111001;
REG[3186] <= 32'b11111100111101001111110000000001;
REG[3187] <= 32'b11111011111110110000000111111011;
REG[3188] <= 32'b11111010000001011111010111111111;
REG[3189] <= 32'b00000001111111011111100111111111;
REG[3190] <= 32'b11110111000001010000010100000011;
REG[3191] <= 32'b00000011000000011111101000001001;
REG[3192] <= 32'b00000110000011010000101011111011;
REG[3193] <= 32'b11110110000001011111010111111000;
REG[3194] <= 32'b00000010000010101111110011111101;
REG[3195] <= 32'b11110011111100100000000000000011;
REG[3196] <= 32'b11111111111111110000001011111101;
REG[3197] <= 32'b00000010000000001111111100001001;
REG[3198] <= 32'b00000010000000000000000011110111;
REG[3199] <= 32'b11110110111101010000110000000000;
REG[3200] <= 32'b11111011111110101111110011110101;
REG[3201] <= 32'b11111111000001101111101111111011;
REG[3202] <= 32'b00000001111101111111101100001011;
REG[3203] <= 32'b00010000111111100000011011110010;
REG[3204] <= 32'b11110100111110111111111011111101;
REG[3205] <= 32'b11111111111110011111111100000001;
REG[3206] <= 32'b00001011000000111111101011111001;
REG[3207] <= 32'b11110011000000011111111000000010;
REG[3208] <= 32'b11111001111101000000000000010111;
REG[3209] <= 32'b00010111000010010000100111111011;
REG[3210] <= 32'b00000010000011000000110100010101;
REG[3211] <= 32'b00010110111111110000011000000110;
REG[3212] <= 32'b11111111000011100000000111111001;
REG[3213] <= 32'b00000001111111100000000100001101;
REG[3214] <= 32'b11110111111101100000011011111100;
REG[3215] <= 32'b00000101111110111111111011111111;
REG[3216] <= 32'b11110110000110010000000100010110;
REG[3217] <= 32'b00000110111110011111000000011011;
REG[3218] <= 32'b00000010000100010000011000010110;
REG[3219] <= 32'b00010100000101101111101000001101;
REG[3220] <= 32'b00000001000001100000010000001010;
REG[3221] <= 32'b00000111111101111111110111111110;
REG[3222] <= 32'b00001000000001100000111011111011;
REG[3223] <= 32'b11111111111110000000100000001001;
REG[3224] <= 32'b00010000111110000000000011111101;
REG[3225] <= 32'b11110100000001000001011000000110;
REG[3226] <= 32'b11111011000010011110100111101111;
REG[3227] <= 32'b00010101000110101111100100001101;
REG[3228] <= 32'b11110101111011010000100000000010;
REG[3229] <= 32'b00000110000010110000110100001000;
REG[3230] <= 32'b00000111111111101110111011111000;
REG[3231] <= 32'b00010010000000110000100100001101;
REG[3232] <= 32'b11111000111110110001101000001001;
REG[3233] <= 32'b00000001111110011111011011111011;
REG[3234] <= 32'b11110010111110001111000011111001;
REG[3235] <= 32'b11111110000000000001110011111101;
REG[3236] <= 32'b00000100111101010000101000000100;
REG[3237] <= 32'b00000001111111001111010011101010;
REG[3238] <= 32'b11111101111111001111001011111100;
REG[3239] <= 32'b00001110111110001111111011111111;
REG[3240] <= 32'b11110010111111110001111000001000;
REG[3241] <= 32'b11111011111111111110111011110111;
REG[3242] <= 32'b00010011000010001111101011111010;
REG[3243] <= 32'b11111001000000010000010100000110;
REG[3244] <= 32'b00000101111110011111100111111110;
REG[3245] <= 32'b00000010000010100001001011111000;
REG[3246] <= 32'b00000110000100100011000111111110;
REG[3247] <= 32'b11111111111111010000110000001110;
REG[3248] <= 32'b00011000111111111111101111111111;
REG[3249] <= 32'b00001110000101100010000111111111;
REG[3250] <= 32'b11110101111110100000010011111100;
REG[3251] <= 32'b00001011111110101111001111111011;
REG[3252] <= 32'b00000001111100010000000011110010;
REG[3253] <= 32'b11110110000010101111001111110010;
REG[3254] <= 32'b11110011111011101111011000001000;
REG[3255] <= 32'b00010010000001110000110000001010;
REG[3256] <= 32'b00001000000001101111100111111100;
REG[3257] <= 32'b11111001111111011111001100000000;
REG[3258] <= 32'b11101101111111011111111011111000;
REG[3259] <= 32'b11101111000000101111111100000101;
REG[3260] <= 32'b11110111111111001111011100000000;
REG[3261] <= 32'b00001001000000000000000000000101;
REG[3262] <= 32'b00000101000000000000101111111011;
REG[3263] <= 32'b11101101111110011111110011111111;
REG[3264] <= 32'b00001001000000001110110100000100;
REG[3265] <= 32'b00001011000001011111100011111100;
REG[3266] <= 32'b11111100111011111111110111111101;
REG[3267] <= 32'b11011110111010111111100011110111;
REG[3268] <= 32'b11110101111111001110001011101010;
REG[3269] <= 32'b11110101111101001111101100000101;
REG[3270] <= 32'b11111101000010011111011111111110;
REG[3271] <= 32'b00001001111101101111010000001110;
REG[3272] <= 32'b00001101111110100000001011101000;
REG[3273] <= 32'b11110001111110111111110011111010;
REG[3274] <= 32'b11110100111101001111101100001001;
REG[3275] <= 32'b00000110111101010000101100001000;
REG[3276] <= 32'b11110100000001000000111011111001;
REG[3277] <= 32'b00000101000001111111010111111011;
REG[3278] <= 32'b00001000111110101111101011110101;
REG[3279] <= 32'b00000011000000111111101111111110;
REG[3280] <= 32'b00000110000010001111110000001101;
REG[3281] <= 32'b00000001000100000000111100010001;
REG[3282] <= 32'b00000000000010000000000100000010;
REG[3283] <= 32'b00000111000000111111111011111111;
REG[3284] <= 32'b11111011111111100000011100001110;
REG[3285] <= 32'b11111110000001101111110000000101;
REG[3286] <= 32'b00000000000010011111101011111110;
REG[3287] <= 32'b11111000000011010000011100001001;
REG[3288] <= 32'b11110110111110011111011011111010;
REG[3289] <= 32'b11110110111101111111101000000010;
REG[3290] <= 32'b00000000000011100000011100000110;
REG[3291] <= 32'b11111100111111110000000100000100;
REG[3292] <= 32'b11110111000000000000011000010101;
REG[3293] <= 32'b11111010111111101111010111111010;
REG[3294] <= 32'b11111110000001111111100100000001;
REG[3295] <= 32'b11111110000001000000000000000001;
REG[3296] <= 32'b11111001111101010000000100001000;
REG[3297] <= 32'b00000110000001101111000111101101;
REG[3298] <= 32'b11110011000000101111011000000011;
REG[3299] <= 32'b11110111111001111111010111110111;
REG[3300] <= 32'b11111011000000001111010011101101;
REG[3301] <= 32'b11111000000001100001101111111110;
REG[3302] <= 32'b11110111000000100000010100000001;
REG[3303] <= 32'b00000000111011101111010011111100;
REG[3304] <= 32'b00000110111111011111110011110111;
REG[3305] <= 32'b11110110111110000000010100000000;
REG[3306] <= 32'b00000110000000101111100111111001;
REG[3307] <= 32'b11101011111101000000000111111101;
REG[3308] <= 32'b00000101111010111101100011101011;
REG[3309] <= 32'b11110110111101001110110011110001;
REG[3310] <= 32'b11100111111101100000001111111011;
REG[3311] <= 32'b11111001111110100000000100000010;
REG[3312] <= 32'b11111110111111011111010111111110;
REG[3313] <= 32'b00000101000000100000001100000010;
REG[3314] <= 32'b11111010000001110000100000000001;
REG[3315] <= 32'b00001100000001101111110111111010;
REG[3316] <= 32'b00000101000000000001011100001010;
REG[3317] <= 32'b00000011000000010000101000000011;
REG[3318] <= 32'b00000101000001010000010000000001;
REG[3319] <= 32'b11110011111111110000110100000111;
REG[3320] <= 32'b11110110111111100000011000000001;
REG[3321] <= 32'b00010011000011011111100011111101;
REG[3322] <= 32'b00000100000010110000011100001000;
REG[3323] <= 32'b11111101111101110000000000000010;
REG[3324] <= 32'b11111110111101000000000011111100;
REG[3325] <= 32'b00001011000000111111110111111110;
REG[3326] <= 32'b11100101000000110000110100001110;
REG[3327] <= 32'b11110001111111101110110111110001;
REG[3328] <= 32'b00000001000011001111001111111011;
REG[3329] <= 32'b11111101111101000000010100000000;
REG[3330] <= 32'b11110010111110111111100111110000;
REG[3331] <= 32'b00000110111110101110100111111010;
REG[3332] <= 32'b11111100111011010000000111111000;
REG[3333] <= 32'b11111010000001100001001000000010;
REG[3334] <= 32'b00000000111111001111001111110000;
REG[3335] <= 32'b11111000111101100000000011111010;
REG[3336] <= 32'b11110001111100111111001011110010;
REG[3337] <= 32'b00000011111110111111011111111010;
REG[3338] <= 32'b11111100000001100000011000000001;
REG[3339] <= 32'b11111000000000011111111000000010;
REG[3340] <= 32'b00001011000010001111101011111110;
REG[3341] <= 32'b11111100000010000000111100000010;
REG[3342] <= 32'b11110100000001011110100111111101;
REG[3343] <= 32'b11111000000000110001001100000101;
REG[3344] <= 32'b11100011000010100000000000000011;
REG[3345] <= 32'b00010100000101011101110111111001;
REG[3346] <= 32'b11110011000000101111000011110011;
REG[3347] <= 32'b11111001000000100000000100000010;
REG[3348] <= 32'b11110011111011011111010100000100;
REG[3349] <= 32'b00001101000000111110111111101011;
REG[3350] <= 32'b11101011000010000000001000000001;
REG[3351] <= 32'b11110111111110110000000100000000;
REG[3352] <= 32'b00000011111111100000001000000101;
REG[3353] <= 32'b00000011000100100001111011111101;
REG[3354] <= 32'b11111001000001010000001000001011;
REG[3355] <= 32'b00001110111101110000000000001101;
REG[3356] <= 32'b00001001111101100000011000001000;
REG[3357] <= 32'b11110110111111000000111011111100;
REG[3358] <= 32'b00000011000010011110101111110100;
REG[3359] <= 32'b00001011000000110000001000001010;
REG[3360] <= 32'b11110010000000011111010011111001;
REG[3361] <= 32'b11111000111101111111100100000001;
REG[3362] <= 32'b11110100111110011111001111110110;
REG[3363] <= 32'b11111111000110011111110100000110;
REG[3364] <= 32'b11111100111111010000111011110010;
REG[3365] <= 32'b11111011111100111111011011111110;
REG[3366] <= 32'b00001110111011111111011111111101;
REG[3367] <= 32'b00000100111111000000000011111001;
REG[3368] <= 32'b00000010111111011111101011110011;
REG[3369] <= 32'b00000100000011010000100000000011;
REG[3370] <= 32'b00000000000000001111010111110111;
REG[3371] <= 32'b11110010111111001111101111110111;
REG[3372] <= 32'b11111001111101011111011000000010;
REG[3373] <= 32'b00010000111111000001000000001100;
REG[3374] <= 32'b00000011111100101110101000000001;
REG[3375] <= 32'b11111011000000110000001000011011;
REG[3376] <= 32'b11110011000001111111011000000010;
REG[3377] <= 32'b00000110111101101111001100000001;
REG[3378] <= 32'b00001000000011000000110100000101;
REG[3379] <= 32'b00000001000010011111011011110111;
REG[3380] <= 32'b11110111000011010000011000001111;
REG[3381] <= 32'b11111000000000101111101000010000;
REG[3382] <= 32'b00000011000010100000001100001100;
REG[3383] <= 32'b00000011000001111111111111111100;
REG[3384] <= 32'b00000001111111101111100100000000;
REG[3385] <= 32'b11110101000000100001000100001011;
REG[3386] <= 32'b00001011111110001111111000001101;
REG[3387] <= 32'b11101100111100011111010100001000;
REG[3388] <= 32'b00010001111110011111010111111100;
REG[3389] <= 32'b11111011000010110001001111111011;
REG[3390] <= 32'b11111100000010000000001000001001;
REG[3391] <= 32'b11110110111011110000011100010110;
REG[3392] <= 32'b00010100000110100001110100011110;
REG[3393] <= 32'b11111000000000001111111100011101;
REG[3394] <= 32'b00010100000011011111001011111000;
REG[3395] <= 32'b11101111000011100000101100001100;
REG[3396] <= 32'b00000000000100011111110111110101;
REG[3397] <= 32'b11111001000001001111010100000101;
REG[3398] <= 32'b00000011111101110000010111111110;
REG[3399] <= 32'b11101111111110000000000000001111;
REG[3400] <= 32'b00010100111011011111010111110001;
REG[3401] <= 32'b11100111000001101110111011111110;
REG[3402] <= 32'b00001010000010011111000000011100;
REG[3403] <= 32'b00000000111101110000010011110101;
REG[3404] <= 32'b11111110000001010000000111110011;
REG[3405] <= 32'b00001100000011100000101000000111;
REG[3406] <= 32'b11111110000000000000111100001101;
REG[3407] <= 32'b00000100000010001111010000000100;
REG[3408] <= 32'b11111000111111111111000000000101;
REG[3409] <= 32'b11110110000001110001001111111100;
REG[3410] <= 32'b11110001111001111110101111111011;
REG[3411] <= 32'b00010101111111011111101111111111;
REG[3412] <= 32'b11111111111110011111010111110101;
REG[3413] <= 32'b00001010000010001111011011111001;
REG[3414] <= 32'b11111000000000111111010100000001;
REG[3415] <= 32'b00100000000010101111001100100110;
REG[3416] <= 32'b11101111111110100000100100001010;
REG[3417] <= 32'b11110101000100001111000111110101;
REG[3418] <= 32'b11111011000000010000011111111110;
REG[3419] <= 32'b00010101111101011111010111111111;
REG[3420] <= 32'b00000110000001010001010011111110;
REG[3421] <= 32'b11111000111111001111111100000000;
REG[3422] <= 32'b00001110111110001111001011111010;
REG[3423] <= 32'b00001101000011100000100100000000;
REG[3424] <= 32'b00000000000011110000001100000100;
REG[3425] <= 32'b00000100111101100000010100001110;
REG[3426] <= 32'b11110111111110100000010000001100;
REG[3427] <= 32'b00000111000010111111100011111011;
REG[3428] <= 32'b00000110111100111111101100001010;
REG[3429] <= 32'b00000110000000000000110111110100;
REG[3430] <= 32'b11110010000001110000100100001000;
REG[3431] <= 32'b00001111111110001111001111111111;
REG[3432] <= 32'b00001111000101000000100000001001;
REG[3433] <= 32'b00001011111100110000000000001010;
REG[3434] <= 32'b00001011000100100000110011110101;
REG[3435] <= 32'b11110100000000111111101000000110;
REG[3436] <= 32'b00001100111110011111101111111101;
REG[3437] <= 32'b00000001000010010000010011111001;
REG[3438] <= 32'b00000001111101001111000000100101;
REG[3439] <= 32'b00001100111110111111111111110111;
REG[3440] <= 32'b00000101000001000000001011110110;
REG[3441] <= 32'b00001110000011100000111111110010;
REG[3442] <= 32'b00000100000000110000100100010111;
REG[3443] <= 32'b00010011111101110000000100000011;
REG[3444] <= 32'b00000001000000010000000011110100;
REG[3445] <= 32'b00000001000000100000000111111011;
REG[3446] <= 32'b11110101111100101111001011110100;
REG[3447] <= 32'b11101111111010111110101000000011;
REG[3448] <= 32'b11101011111100101111000111111001;
REG[3449] <= 32'b11110001000010001111000111101010;
REG[3450] <= 32'b00000111000000111111111100001100;
REG[3451] <= 32'b00000110000000110000011000000001;
REG[3452] <= 32'b11110011000001011111111011111001;
REG[3453] <= 32'b00010000000100100000000111111110;
REG[3454] <= 32'b11111101111110111111111111111010;
REG[3455] <= 32'b11111011111111101111101011111000;
REG[3456] <= 32'b00000101000001110000101111111001;
REG[3457] <= 32'b11110011111111011111011011111111;
REG[3458] <= 32'b11111011000001101111110011111001;
REG[3459] <= 32'b00010111000001110000010000000110;
REG[3460] <= 32'b00001001111110100000011011110111;
REG[3461] <= 32'b00000011000000100000010111111110;
REG[3462] <= 32'b00100101111110100000000111111010;
REG[3463] <= 32'b11111001111110101111010100000101;
REG[3464] <= 32'b11111110111010001111111000010101;
REG[3465] <= 32'b11111101000001001111111011110011;
REG[3466] <= 32'b11111001111110001111110011110111;
REG[3467] <= 32'b11110110111101000000001111111011;
REG[3468] <= 32'b11110111000001001111101100000010;
REG[3469] <= 32'b00001010111111001111110100000000;
REG[3470] <= 32'b11111111111111100000100111110010;
REG[3471] <= 32'b00001110111111011111101100000101;
REG[3472] <= 32'b00000101111111000000010111110111;
REG[3473] <= 32'b11111100000001000001001100001101;
REG[3474] <= 32'b00001010111100111111001000000101;
REG[3475] <= 32'b11110101111110010000011100000000;
REG[3476] <= 32'b11111001000000000000011011111100;
REG[3477] <= 32'b00000011000000010001101111110010;
REG[3478] <= 32'b00000011000010101111010111111010;
REG[3479] <= 32'b00010001111110000000001100001010;
REG[3480] <= 32'b11110001111100110000001111110010;
REG[3481] <= 32'b11110100111111010000011000001011;
REG[3482] <= 32'b00000101111001101111000000000110;
REG[3483] <= 32'b00001001111111010000001111110001;
REG[3484] <= 32'b11101110111111100000011100000101;
REG[3485] <= 32'b00000001111110011111001011111110;
REG[3486] <= 32'b00000101000011100001000011111010;
REG[3487] <= 32'b11111101000001111111101011111011;
REG[3488] <= 32'b00000011111110001111101111111111;
REG[3489] <= 32'b11111011111010011110101011111000;
REG[3490] <= 32'b11111001111111101110110000000101;
REG[3491] <= 32'b11101100000000110000101011111111;
REG[3492] <= 32'b11101100111111111111001111111110;
REG[3493] <= 32'b11111101000000011111000000001001;
REG[3494] <= 32'b11110010000000010000000111111111;
REG[3495] <= 32'b00010110000011100001000100000000;
REG[3496] <= 32'b00000101000000010000000111111010;
REG[3497] <= 32'b11110111000001110000100000000010;
REG[3498] <= 32'b11110111111111011111101011111110;
REG[3499] <= 32'b00000001111111100000100000000001;
REG[3500] <= 32'b00000000111101111111110000001111;
REG[3501] <= 32'b00000001111110001111101011101100;
REG[3502] <= 32'b11101110000101000000111000001001;
REG[3503] <= 32'b11111110111101111111011100001001;
REG[3504] <= 32'b11110000111110010000000111111000;
REG[3505] <= 32'b00000001000000001111100000000000;
REG[3506] <= 32'b00001100000010100001000100001000;
REG[3507] <= 32'b11101010000000110001110100000000;
REG[3508] <= 32'b00000110000010111111010111110110;
REG[3509] <= 32'b11111100111110110000001011111110;
REG[3510] <= 32'b11111011111110000001010000001001;
REG[3511] <= 32'b00001011000001001111010111101101;
REG[3512] <= 32'b00000100111111010000010111111101;
REG[3513] <= 32'b11101110111010011111110000000111;
REG[3514] <= 32'b11111110000010101111000111011101;
REG[3515] <= 32'b11101011000101100000011011111110;
REG[3516] <= 32'b00010111111101011111001111110010;
REG[3517] <= 32'b00001011000010101111010000001010;
REG[3518] <= 32'b11101011111010101110000011110101;
REG[3519] <= 32'b00000101011100100000001011101000;
REG[3520] <= 32'b11110000111101111111100100000010;
REG[3521] <= 32'b11100011111100111111101111111110;
REG[3522] <= 32'b11101110111110111111111100001010;
REG[3523] <= 32'b11111101000001111110101111111011;
REG[3524] <= 32'b00000001000000011111100011111001;
REG[3525] <= 32'b11110001111101001111010000000100;
REG[3526] <= 32'b00000010000000001111100011111000;
REG[3527] <= 32'b11111011111110101111010111110011;
REG[3528] <= 32'b00000101111110010000011011111101;
REG[3529] <= 32'b11110100111110001111111111110111;
REG[3530] <= 32'b00000001111111101111100011110110;
REG[3531] <= 32'b11110101111110001111100111111110;
REG[3532] <= 32'b00001011000010111111010111111011;
REG[3533] <= 32'b00000000000011000000111100001111;
REG[3534] <= 32'b11111001111101011111101000000010;
REG[3535] <= 32'b11111101111100101111110111111100;
REG[3536] <= 32'b11111100000001110000011100000011;
REG[3537] <= 32'b11111101111110001111110011110111;
REG[3538] <= 32'b11111110111110010000000111111000;
REG[3539] <= 32'b11110111000010110001100000001000;
REG[3540] <= 32'b11111010111111000001100011110111;
REG[3541] <= 32'b00011100111010110000101000000001;
REG[3542] <= 32'b00001000000001000010100111101010;
REG[3543] <= 32'b00001101000001100000011011100001;
REG[3544] <= 32'b11101111111100000001111100000101;
REG[3545] <= 32'b11110011111111101111110111111010;
REG[3546] <= 32'b00011101111110011110101100000001;
REG[3547] <= 32'b00000001111110100000010111111100;
REG[3548] <= 32'b11111101000001111111110011111100;
REG[3549] <= 32'b11111110111110011111110000000100;
REG[3550] <= 32'b11111000111111010000111100001101;
REG[3551] <= 32'b00000010000011000011101000001101;
REG[3552] <= 32'b00001001000001000000001011111000;
REG[3553] <= 32'b00010110000101000000000011110000;
REG[3554] <= 32'b11110001000001001111011011110110;
REG[3555] <= 32'b11111011111101000001000000000010;
REG[3556] <= 32'b00001110000000111111111011110111;
REG[3557] <= 32'b00001000000010000001011100001000;
REG[3558] <= 32'b11111001000000111111111100001111;
REG[3559] <= 32'b11110001111011101111011000000111;
REG[3560] <= 32'b00000100000011011111010111101100;
REG[3561] <= 32'b11101110000000000000000000010010;
REG[3562] <= 32'b11111000111101000001001100000011;
REG[3563] <= 32'b11110110111110010000101100001010;
REG[3564] <= 32'b00001001111100101111001000000010;
REG[3565] <= 32'b00010011000100010000100100001000;
REG[3566] <= 32'b11111100111110001111111100001100;
REG[3567] <= 32'b00000010111101111110111100000100;
REG[3568] <= 32'b11111100000000101111010111110110;
REG[3569] <= 32'b11110010111110001111101011111110;
REG[3570] <= 32'b11110101111101111111101011111110;
REG[3571] <= 32'b00001001000001111111111111110101;
REG[3572] <= 32'b11101101111101001111010011111010;
REG[3573] <= 32'b00000011111100001110110111101101;
REG[3574] <= 32'b11101110111101100000101011101000;
REG[3575] <= 32'b11110001111101011111100011110010;
REG[3576] <= 32'b11111011000001111111100000001110;
REG[3577] <= 32'b00001011111100001111110011111001;
REG[3578] <= 32'b11111101000001110000010011111000;
REG[3579] <= 32'b11111111111111100001000111111010;
REG[3580] <= 32'b11110111111011111111011111110011;
REG[3581] <= 32'b11111000001000100000111111101010;
REG[3582] <= 32'b00000001111100100000010100010011;
REG[3583] <= 32'b00100101111101010000000111110011;
REG[3584] <= 32'b00000001000001000001110011111111;
REG[3585] <= 32'b11111001111111000000000000011111;
REG[3586] <= 32'b00000011111100100000100000001000;
REG[3587] <= 32'b11111101000110010000111111101100;
REG[3588] <= 32'b00010000000011111111111100001100;
REG[3589] <= 32'b11111100111100001110110111110110;
REG[3590] <= 32'b00000011000000011111111100000111;
REG[3591] <= 32'b11111011000010101111111100000101;
REG[3592] <= 32'b11111001000000011111011100010011;
REG[3593] <= 32'b00010001000011001111101011111010;
REG[3594] <= 32'b11100101000000000000100111110111;
REG[3595] <= 32'b00000101000111000011000100100011;
REG[3596] <= 32'b00000100111111010001000100100011;
REG[3597] <= 32'b00000001000010001111001000000001;
REG[3598] <= 32'b00000000000010011111011111111100;
REG[3599] <= 32'b11110100000010000000011011111100;
REG[3600] <= 32'b11110101111101111110111100001000;
REG[3601] <= 32'b00000110111111011111001111110111;
REG[3602] <= 32'b11110101111110010000000011111011;
REG[3603] <= 32'b00001100000001000000001011110111;
REG[3604] <= 32'b00000100000000100000011000000101;
REG[3605] <= 32'b00000101111100111111111111111111;
REG[3606] <= 32'b00001010111101001111010011111001;
REG[3607] <= 32'b11110000111110111111001111111000;
REG[3608] <= 32'b00000111000011100000110100001000;
REG[3609] <= 32'b11111011111110100000101000000001;
REG[3610] <= 32'b00000101111111001111111111110101;
REG[3611] <= 32'b00001101000000000001011100001101;
REG[3612] <= 32'b00000000111011101111001000001100;
REG[3613] <= 32'b00010010000000100000001011111001;
REG[3614] <= 32'b00001110000000101111110111111001;
REG[3615] <= 32'b00001111000010010001001100000110;
REG[3616] <= 32'b00000111111111000001000111111010;
REG[3617] <= 32'b11110001111011101111000011111001;
REG[3618] <= 32'b00010001111000111110101111111010;
REG[3619] <= 32'b00000100000001100010010100010010;
REG[3620] <= 32'b11011000000000000000111000000101;
REG[3621] <= 32'b00000011111110001111101011111011;
REG[3622] <= 32'b00000000000001101111111111110110;
REG[3623] <= 32'b11110010000000010000100011111000;
REG[3624] <= 32'b11111011111010111110101111111111;
REG[3625] <= 32'b11111101111111111111110000010000;
REG[3626] <= 32'b00001010000000000000101000000010;
REG[3627] <= 32'b11110110111111110000100000000010;
REG[3628] <= 32'b00010101111111001111111000000101;
REG[3629] <= 32'b00100010000010100010010111111100;
REG[3630] <= 32'b11111110000001011111101011111010;
REG[3631] <= 32'b11111000000010001111000111111110;
REG[3632] <= 32'b11110010111111101111110011111101;
REG[3633] <= 32'b11111011111110101111011011111011;
REG[3634] <= 32'b11110101000001101111001011110110;
REG[3635] <= 32'b11111001111101111111100100000010;
REG[3636] <= 32'b00011101010010000001110011110110;
REG[3637] <= 32'b11110110111101110000111000100010;
REG[3638] <= 32'b00011000111110111111101111111100;
REG[3639] <= 32'b00000000111111001111101111111101;
REG[3640] <= 32'b11111010111111111111100111110110;
REG[3641] <= 32'b11110111111111010000100100000011;
REG[3642] <= 32'b11110110111110001111111000000001;
REG[3643] <= 32'b00001010000001111111010011110010;
REG[3644] <= 32'b11110110111111011111101011111010;
REG[3645] <= 32'b00001000111111001111110111111011;
REG[3646] <= 32'b11111000111111010000011011111100;
REG[3647] <= 32'b11111101111100111111001100000010;
REG[3648] <= 32'b11111110111101011111110100010100;
REG[3649] <= 32'b00010000000011111111111011110011;
REG[3650] <= 32'b11111111000100000001000000011000;
REG[3651] <= 32'b11111000111010111111010100001111;
REG[3652] <= 32'b00001001000011001111100100000110;
REG[3653] <= 32'b00001001111111111111110011111010;
REG[3654] <= 32'b11110101111111110000011111111110;
REG[3655] <= 32'b11111100111111010000001100001101;
REG[3656] <= 32'b00001011111110101111100111111010;
REG[3657] <= 32'b00000010111110001111111111111111;
REG[3658] <= 32'b11111000000000100000001011110000;
REG[3659] <= 32'b11111100111111101111101011111110;
REG[3660] <= 32'b11111110111111000000010011111100;
REG[3661] <= 32'b11110011000001010000011000011000;
REG[3662] <= 32'b00001010000000000000001011110110;
REG[3663] <= 32'b11101010111100101111001100000011;
REG[3664] <= 32'b00000011111101001111010100000000;
REG[3665] <= 32'b00000101000001010000100011111010;
REG[3666] <= 32'b11111101000000010000011011111000;
REG[3667] <= 32'b11110011111101110000000000000010;
REG[3668] <= 32'b00000111111110011111001011111001;
REG[3669] <= 32'b11111111000000001111110011111011;
REG[3670] <= 32'b11110100111101000000111100001101;
REG[3671] <= 32'b00000010000000101111111011111110;
REG[3672] <= 32'b11111100111010101110111000000010;
REG[3673] <= 32'b11111010000000111111011111110111;
REG[3674] <= 32'b11111100111111111111100100000001;
REG[3675] <= 32'b11101110111110001111001100000010;
REG[3676] <= 32'b11111010111110000000110100011101;
REG[3677] <= 32'b00000011000001010000000011111010;
REG[3678] <= 32'b11101010111101111110111011111110;
REG[3679] <= 32'b11111011111101010000000111110110;
REG[3680] <= 32'b11110001111111010000000111111110;
REG[3681] <= 32'b11111001111101011111100100000010;
REG[3682] <= 32'b00000101111110110000001111111101;
REG[3683] <= 32'b11110100000000100000000111110101;
REG[3684] <= 32'b11110110111110110000010011101111;
REG[3685] <= 32'b11110100111111111111101011111101;
REG[3686] <= 32'b00001010111001101111010111110111;
REG[3687] <= 32'b00000000000000000000011011101101;
REG[3688] <= 32'b11110100000010100001011000000100;
REG[3689] <= 32'b11110101000001010000000100001000;
REG[3690] <= 32'b11101101111101010000001011111101;
REG[3691] <= 32'b11111010000001111111101000000001;
REG[3692] <= 32'b11111011111111101111111100000111;
REG[3693] <= 32'b00000000000000111111111100000000;
REG[3694] <= 32'b11111101111111101111100111111111;
REG[3695] <= 32'b11110111111100110000010011111000;
REG[3696] <= 32'b11110110000000011111110011110110;
REG[3697] <= 32'b00001000000001000010011100010001;
REG[3698] <= 32'b00010110000000000000001100000111;
REG[3699] <= 32'b11110111111011001111100111111101;
REG[3700] <= 32'b11111110000000111111010111111110;
REG[3701] <= 32'b11111111111111110000010100000011;
REG[3702] <= 32'b11110011111111010000010100000100;
REG[3703] <= 32'b00000010111111111111000000000000;
REG[3704] <= 32'b00000010000001100000001100001000;
REG[3705] <= 32'b11110100000000000000001011110110;
REG[3706] <= 32'b11111001111111010000100111110000;
REG[3707] <= 32'b11110111111111001111010011111010;
REG[3708] <= 32'b00001000111111011111010011111011;
REG[3709] <= 32'b11110111111111110000101000000110;
REG[3710] <= 32'b11111111000001101111101100000001;
REG[3711] <= 32'b00010001000010010001011111111110;
REG[3712] <= 32'b00001000000001000010010000011000;
REG[3713] <= 32'b00100011111111100000010000000100;
REG[3714] <= 32'b00100001000101110010100000000011;
REG[3715] <= 32'b00000010000001011111100011101010;
REG[3716] <= 32'b11110101111101101111101100000111;
REG[3717] <= 32'b11110001111010110000100111111101;
REG[3718] <= 32'b00000110000011110000010000000111;
REG[3719] <= 32'b00010000111110111111111100000101;
REG[3720] <= 32'b11111100111111100000000111111111;
REG[3721] <= 32'b11111110111101111111111000000011;
REG[3722] <= 32'b00001000000000011111110011110111;
REG[3723] <= 32'b11111000111110110000010000001101;
REG[3724] <= 32'b11111111111010100011000000011001;
REG[3725] <= 32'b00001011111101011111111111100010;
REG[3726] <= 32'b11111010111111010000001100000100;
REG[3727] <= 32'b00100100111100100000100100010001;
REG[3728] <= 32'b00000011111111000001000011101111;
REG[3729] <= 32'b00000001000001001111110100001010;
REG[3730] <= 32'b11111110111111011111110000000101;
REG[3731] <= 32'b11111100000001001111110111111100;
REG[3732] <= 32'b00000011000001010000001000000010;
REG[3733] <= 32'b11110111111111100000010100000110;
REG[3734] <= 32'b11111101111111111111111000001010;
REG[3735] <= 32'b11110100000010011111010011111110;
REG[3736] <= 32'b11111100000010010000000100000110;
REG[3737] <= 32'b11110100111111110000000000001011;
REG[3738] <= 32'b11110110111111101111101011101000;
REG[3739] <= 32'b11111001111110011111111000001000;
REG[3740] <= 32'b00000000111001110000000111111011;
REG[3741] <= 32'b11111111000000101111110111101000;
REG[3742] <= 32'b11110101111111011111111000000011;
REG[3743] <= 32'b11101110000001010000000011111100;
REG[3744] <= 32'b00000100000000111111010011111110;
REG[3745] <= 32'b11111101111111110000011000000100;
REG[3746] <= 32'b00001000000000101111110000000000;
REG[3747] <= 32'b11110100111111010000000100000100;
REG[3748] <= 32'b00000011000000111111111100001000;
REG[3749] <= 32'b00010100000010100000101000010010;
REG[3750] <= 32'b11111110111110000000001000010011;
REG[3751] <= 32'b00000110000010111111101011110111;
REG[3752] <= 32'b11110001111101001111111011111000;
REG[3753] <= 32'b11110011111010011111011011110100;
REG[3754] <= 32'b11111110111101101111111011110011;
REG[3755] <= 32'b11111111111100100000000011111100;
REG[3756] <= 32'b11101010111101001111101111111000;
REG[3757] <= 32'b11110011111101111111101011111010;
REG[3758] <= 32'b00000001111100001110011111111111;
REG[3759] <= 32'b00000000000000000000001011110110;
REG[3760] <= 32'b11110111000000001111001011110000;
REG[3761] <= 32'b11110011111101001111100000000101;
REG[3762] <= 32'b11110000111110001111100111101110;
REG[3763] <= 32'b00000000000011011111101011110011;
REG[3764] <= 32'b11111001111100111111110100000010;
REG[3765] <= 32'b11111000111100111111101011111000;
REG[3766] <= 32'b11110110111101011111011011111001;
REG[3767] <= 32'b00000001111111001111100100000100;
REG[3768] <= 32'b11111110000000011111111100000101;
REG[3769] <= 32'b11111010111111100000001011110010;
REG[3770] <= 32'b00000110111101010000001111111011;
REG[3771] <= 32'b11101011111100001111011111110001;
REG[3772] <= 32'b00000101111101011111001111111001;
REG[3773] <= 32'b11110111111110110000011011110100;
REG[3774] <= 32'b00000011000010000000100100000111;
REG[3775] <= 32'b00000000111111011111110100000100;
REG[3776] <= 32'b00000011000010111111111111110111;
REG[3777] <= 32'b11111111000000110000101100001001;
REG[3778] <= 32'b00000100000000111111100111101001;
REG[3779] <= 32'b11111010111111111111101000001111;
REG[3780] <= 32'b00000100111101011111010011110010;
REG[3781] <= 32'b11101110000010110001110000000111;
REG[3782] <= 32'b11111111111111011111110100010001;
REG[3783] <= 32'b11111111000110010001001100000100;
REG[3784] <= 32'b11111111000010111111011100001011;
REG[3785] <= 32'b00001001111111001111100100000101;
REG[3786] <= 32'b11111110000010110000111000000100;
REG[3787] <= 32'b00000010000001100000111011111100;
REG[3788] <= 32'b11110111000001001111011111111010;
REG[3789] <= 32'b00001000000010111111111000000101;
REG[3790] <= 32'b11110110111111100000100000100011;
REG[3791] <= 32'b00010101000011001111111100000101;
REG[3792] <= 32'b11111001111101101111101111111101;
REG[3793] <= 32'b11110011111010111110110011100111;
REG[3794] <= 32'b11110110111110101110111111100111;
REG[3795] <= 32'b11110011111011101111011011111111;
REG[3796] <= 32'b11111000111110000000100111111010;
REG[3797] <= 32'b11111010111101011111011111111000;
REG[3798] <= 32'b00000110111110011111000111111110;
REG[3799] <= 32'b00001010111111110000000000000011;
REG[3800] <= 32'b11111000000000100000011011101101;
REG[3801] <= 32'b00001000111110111111110111111101;
REG[3802] <= 32'b11111111000010010000111111110111;
REG[3803] <= 32'b11111101000001100001001000001011;
REG[3804] <= 32'b00000000111111011111110111111100;
REG[3805] <= 32'b00000101000011001111100111101110;
REG[3806] <= 32'b11111110000100000000011000010110;
REG[3807] <= 32'b00000100111110010000011000000010;
REG[3808] <= 32'b00001000000010011111110111111000;
REG[3809] <= 32'b11110111000100000001111011111000;
REG[3810] <= 32'b00001011000100010000110111111100;
REG[3811] <= 32'b00000000111111000000001100000000;
REG[3812] <= 32'b00001001111101101111010011111001;
REG[3813] <= 32'b11110011111100100000011111111011;
REG[3814] <= 32'b11110111000001100000011000010001;
REG[3815] <= 32'b00000100111111011111100111111101;
REG[3816] <= 32'b00010000000010101111111011111011;
REG[3817] <= 32'b11111100000011000001001000000111;
REG[3818] <= 32'b00001000111111010000101100001001;
REG[3819] <= 32'b00001100111110010000101111111100;
REG[3820] <= 32'b11111010111110110000101111110111;
REG[3821] <= 32'b00000011000001011111110100000011;
REG[3822] <= 32'b11111110111101101111110111111101;
REG[3823] <= 32'b11110100000001000000010000001010;
REG[3824] <= 32'b11111110000010010000010100001010;
REG[3825] <= 32'b11110111111111100000000100001100;
REG[3826] <= 32'b11111111000000011111110011111101;
REG[3827] <= 32'b11111011111100001110101011110011;
REG[3828] <= 32'b00000010111101001111111111111110;
REG[3829] <= 32'b11111010000000011111011100000101;
REG[3830] <= 32'b11111111111110111110111000000011;
REG[3831] <= 32'b11110010111101010000000100001010;
REG[3832] <= 32'b00000011000011110000001111110011;
REG[3833] <= 32'b11111010111111001111011100000011;
REG[3834] <= 32'b00001110111111001111011100001100;
REG[3835] <= 32'b11111011000011001110101111110010;
REG[3836] <= 32'b11111110111110110000100100001100;
REG[3837] <= 32'b00000000000000001111111100000110;
REG[3838] <= 32'b00000010111111011111100100000011;
REG[3839] <= 32'b11111010000001000000000111110111;
REG[3840] <= 32'b00000010000000101111011100000010;
REG[3841] <= 32'b11111111111101001111111111110011;
REG[3842] <= 32'b11111101111110000000011011111110;
REG[3843] <= 32'b00001010111101001111111100010001;
REG[3844] <= 32'b11110010111111101111100111110000;
REG[3845] <= 32'b11111011111101101111100100001010;
REG[3846] <= 32'b00000000111100101111110111111100;
REG[3847] <= 32'b11111000111111011111101111110000;
REG[3848] <= 32'b11111111111101101111000111110100;
REG[3849] <= 32'b11110111111110001111110100000101;
REG[3850] <= 32'b00000101000000011110101111110010;
REG[3851] <= 32'b00001110000001101111010011110111;
REG[3852] <= 32'b11110001111110100000110000000000;
REG[3853] <= 32'b11111101111110101110110111111111;
REG[3854] <= 32'b00011110111110111111111100001001;
REG[3855] <= 32'b00010101000010110000010000000101;
REG[3856] <= 32'b00001100000001010001111000001111;
REG[3857] <= 32'b00000101000110110001100000001100;
REG[3858] <= 32'b00010111000010011111100100010100;
REG[3859] <= 32'b00010001000100010000001111111010;
REG[3860] <= 32'b11110001111011011111011111111100;
REG[3861] <= 32'b00001001000000010000010111110000;
REG[3862] <= 32'b11110011111101110000010011111001;
REG[3863] <= 32'b11110111111110110000001011110110;
REG[3864] <= 32'b00010011111111111111010011110110;
REG[3865] <= 32'b00000110111111001111111011111010;
REG[3866] <= 32'b11110111111110100000111011111110;
REG[3867] <= 32'b00001100111110110000010011110010;
REG[3868] <= 32'b00001000111111010000010100001100;
REG[3869] <= 32'b00000001111111011110100111111100;
REG[3870] <= 32'b00000100000101010000111000000111;
REG[3871] <= 32'b11110100111111111111010000000010;
REG[3872] <= 32'b11111011111101101111101100001000;
REG[3873] <= 32'b00010011111111011111010100000000;
REG[3874] <= 32'b11111000000011000011000111111111;
REG[3875] <= 32'b11111000111101101111000100000000;
REG[3876] <= 32'b00010101111110001111000111110111;
REG[3877] <= 32'b11110100000000111111010100000000;
REG[3878] <= 32'b11111100111111011111011000000111;
REG[3879] <= 32'b00000011000000001111110011111011;
REG[3880] <= 32'b11110011000001000000011011111111;
REG[3881] <= 32'b11111010111011101111011100000000;
REG[3882] <= 32'b11110110111101011110100111111110;
REG[3883] <= 32'b11110101111101101111001111111000;
REG[3884] <= 32'b11101101111110101111001111101110;
REG[3885] <= 32'b11111000000000001111001111111001;
REG[3886] <= 32'b11110101111101111111011011111111;
REG[3887] <= 32'b00001100000010110000000011110100;
REG[3888] <= 32'b11111011111101100000010100000100;
REG[3889] <= 32'b11111100000000111111001111110011;
REG[3890] <= 32'b00000101111101110000010000001000;
REG[3891] <= 32'b11110011111110100000010000000100;
REG[3892] <= 32'b00000010000100001111101011111101;
REG[3893] <= 32'b00000010111111111111010000000101;
REG[3894] <= 32'b11110110111111110001000000000101;
REG[3895] <= 32'b11111111000101111111111011111000;
REG[3896] <= 32'b11110101110111111111001011101100;
REG[3897] <= 32'b00000000111110001111010111101100;
REG[3898] <= 32'b11111000111101001111110011101110;
REG[3899] <= 32'b11110000111111101111110011110110;
REG[3900] <= 32'b00001100111111010000011100000111;
REG[3901] <= 32'b00001011000001101111111000000111;
REG[3902] <= 32'b11111011000001001111001111111010;
REG[3903] <= 32'b11110110000000001111110011111001;
REG[3904] <= 32'b11111101111110100000111000010010;
REG[3905] <= 32'b00000101111111111111100011111111;
REG[3906] <= 32'b11111111000010000000011011111011;
REG[3907] <= 32'b11101110111110111111110100001011;
REG[3908] <= 32'b00000101111111110000000000000100;
REG[3909] <= 32'b11110000111110010000011011111001;
REG[3910] <= 32'b11111110111111101110111111111111;
REG[3911] <= 32'b00010011000001100001001111111111;
REG[3912] <= 32'b11110011000000010001100000000110;
REG[3913] <= 32'b00000110111111010000000011111001;
REG[3914] <= 32'b00010101000000001111001100000001;
REG[3915] <= 32'b11110010111111000001000000010001;
REG[3916] <= 32'b00000001000001011111101100000010;
REG[3917] <= 32'b00101000111110110000001100011000;
REG[3918] <= 32'b11111111111110011111001011111110;
REG[3919] <= 32'b11111111000001111111110111110010;
REG[3920] <= 32'b11101010111110001111100011111111;
REG[3921] <= 32'b11101111000000001111000111111101;
REG[3922] <= 32'b00000000000001101111001111111001;
REG[3923] <= 32'b11110000000010101111110111111101;
REG[3924] <= 32'b11101011111101000000000111111011;
REG[3925] <= 32'b11111100000100011111001111110111;
REG[3926] <= 32'b11101111000000110000110100000101;
REG[3927] <= 32'b00010100000110111110110011111001;
REG[3928] <= 32'b11110011000010100001100100010111;
REG[3929] <= 32'b11111101000101110001000100010110;
REG[3930] <= 32'b00000110111111011110111011111100;
REG[3931] <= 32'b11111000000000100001010100000100;
REG[3932] <= 32'b00000010111110011111110111111001;
REG[3933] <= 32'b00010011000010010000110111110111;
REG[3934] <= 32'b11111101111111110000111100000100;
REG[3935] <= 32'b11111100000000010000000100000101;
REG[3936] <= 32'b11111000111101111111110111101010;
REG[3937] <= 32'b11110000111011011111000011111100;
REG[3938] <= 32'b11111010111011001111000111101110;
REG[3939] <= 32'b11101101111110011111101011101110;
REG[3940] <= 32'b11110001111101000000000000001101;
REG[3941] <= 32'b00101000111111111111111100001010;
REG[3942] <= 32'b00000011000011100000110000001001;
REG[3943] <= 32'b00001111000100000000000111101110;
REG[3944] <= 32'b11110000000000110000111100010111;
REG[3945] <= 32'b00000110111110101111100011111000;
REG[3946] <= 32'b11111110000001010000000011111001;
REG[3947] <= 32'b00000101111100100000011000000100;
REG[3948] <= 32'b11111101111100010000001011111010;
REG[3949] <= 32'b00000101111111000000001111101011;
REG[3950] <= 32'b11110101000001011111100000000100;
REG[3951] <= 32'b11111110111011101111110000010011;
REG[3952] <= 32'b00000101000001011111101011111100;
REG[3953] <= 32'b00000010000010100000000000001110;
REG[3954] <= 32'b00000100000000111111111100000010;
REG[3955] <= 32'b00001000000001100010011000011001;
REG[3956] <= 32'b00000000111111010000101100001010;
REG[3957] <= 32'b00110010000111111111101011111000;
REG[3958] <= 32'b11111100111111101110111011111111;
REG[3959] <= 32'b11110110111110111110111111110011;
REG[3960] <= 32'b00000010111111101110010000000000;
REG[3961] <= 32'b11111010111100000000100111110000;
REG[3962] <= 32'b11100111111111011111100011101111;
REG[3963] <= 32'b11111011000000010000100011111100;
REG[3964] <= 32'b11110101111110001111011111111110;
REG[3965] <= 32'b00000110111111001111100111111101;
REG[3966] <= 32'b11111011111101111111011011111011;
REG[3967] <= 32'b11110010111101001111000111110111;
REG[3968] <= 32'b00000000111011000000010100010010;
REG[3969] <= 32'b11110010111101101111010111110010;
REG[3970] <= 32'b00000000000011101111011111111100;
REG[3971] <= 32'b11111010111110011111111100000110;
REG[3972] <= 32'b11110011111011100000010111111011;
REG[3973] <= 32'b11101000111101101111011011101001;
REG[3974] <= 32'b00000000111101011110000111110011;
REG[3975] <= 32'b00000110000000110000101100100001;
REG[3976] <= 32'b00001001000011011111010100000001;
REG[3977] <= 32'b00011010111011101111010100010101;
REG[3978] <= 32'b11111000111111111111110100000010;
REG[3979] <= 32'b00000011000101001111010011111101;
REG[3980] <= 32'b11110111111010111111011000001100;
REG[3981] <= 32'b11111100111111010000001100000011;
REG[3982] <= 32'b11110010000001111111011011110110;
REG[3983] <= 32'b00000001111100101110101100000101;
REG[3984] <= 32'b11110110111101001111111000001100;
REG[3985] <= 32'b11111011000001001111000111110010;
REG[3986] <= 32'b11100101000000111111010111111000;
REG[3987] <= 32'b11110010111011111110100111111110;
REG[3988] <= 32'b00000100000010001111111011111110;
REG[3989] <= 32'b11111001111100011111011000011000;
REG[3990] <= 32'b11110101111111011111101111110011;
REG[3991] <= 32'b11110101000000111111111011111101;
REG[3992] <= 32'b11111110111101001111011100000000;
REG[3993] <= 32'b00001000111110001111111011111010;
REG[3994] <= 32'b11111100000001000000101100000011;
REG[3995] <= 32'b11110111000010101111101100000000;
REG[3996] <= 32'b00001101001000100000100000001011;
REG[3997] <= 32'b11111100000001000000010100000010;
REG[3998] <= 32'b00000011111111111111011000000010;
REG[3999] <= 32'b00010001111111101111011100010010;
REG[4000] <= 32'b00010110000110000001111000001011;
REG[4001] <= 32'b11101010000100000000100000000000;
REG[4002] <= 32'b00101001001000000000001000001011;
REG[4003] <= 32'b00000001000000001111100011110110;
REG[4004] <= 32'b11111001000000001111110111111000;
REG[4005] <= 32'b11110100111110001111100000000010;
REG[4006] <= 32'b00000110111110111111010011111010;
REG[4007] <= 32'b11110010000001101111111011111100;
REG[4008] <= 32'b11111011111111111111111000000110;
REG[4009] <= 32'b00000100000000001111100111111011;
REG[4010] <= 32'b11111000111110001111011011111101;
REG[4011] <= 32'b11111011111110101111110011111110;
REG[4012] <= 32'b11110101111101111111101100000100;
REG[4013] <= 32'b11111101000000110000011100011101;
REG[4014] <= 32'b00000000000001100000010011111101;
REG[4015] <= 32'b11110000000111001111011000001110;
REG[4016] <= 32'b00001001111111111111101100000001;
REG[4017] <= 32'b11111111000000110000100111110101;
REG[4018] <= 32'b11110011000001001111110100000001;
REG[4019] <= 32'b00000011111011111110111011111011;
REG[4020] <= 32'b11111110111111100000010000000100;
REG[4021] <= 32'b11110110111110000000100000001001;
REG[4022] <= 32'b11111001000010001111100011111001;
REG[4023] <= 32'b00101001001000011111101000010110;
REG[4024] <= 32'b11111101111101100010001100010100;
REG[4025] <= 32'b11111111000101100000000011110101;
REG[4026] <= 32'b00001100000001100000000000001111;
REG[4027] <= 32'b00000011000000110001110000001010;
REG[4028] <= 32'b11111111000001101111101111111001;
REG[4029] <= 32'b00010111000100000000011000000010;
REG[4030] <= 32'b11111110111110001111110000000010;
REG[4031] <= 32'b11111001111011110000101000111100;
REG[4032] <= 32'b00001111000011111111111011110010;
REG[4033] <= 32'b00001011001100110001010100010010;
REG[4034] <= 32'b00000101111011001111011100001101;
REG[4035] <= 32'b11110010111101010000011100100101;
REG[4036] <= 32'b00011111000101001111010111111000;
REG[4037] <= 32'b00000011000100010001000000001110;
REG[4038] <= 32'b11101111111101111111011100010011;
REG[4039] <= 32'b00010111000011010001001100100001;
REG[4040] <= 32'b00011100000000000000010000001101;
REG[4041] <= 32'b00010000000011100001100111111001;
REG[4042] <= 32'b00010000000010000001011100001011;
REG[4043] <= 32'b00010000111100110000001100000110;
REG[4044] <= 32'b11111000000001000000010111111001;
REG[4045] <= 32'b11110100000000101111100000000110;
REG[4046] <= 32'b11111110111100101110110100001011;
REG[4047] <= 32'b11110000111111111111111111110101;
REG[4048] <= 32'b11111000111110111110111111111010;
REG[4049] <= 32'b11111111000000001111111000000010;
REG[4050] <= 32'b11111001111110111111100111110101;
REG[4051] <= 32'b11111011000000001111001111101111;
REG[4052] <= 32'b11101111111110011111010100001101;
REG[4053] <= 32'b11111010000001010001010011111000;
REG[4054] <= 32'b00001011000001001111000011111001;
REG[4055] <= 32'b00001010000000000001101100010000;
REG[4056] <= 32'b11110010111111010000100111111000;
REG[4057] <= 32'b00001000000000101111000011110001;
REG[4058] <= 32'b11110000111110110000000100010111;
REG[4059] <= 32'b11111110111101001111100111110001;
REG[4060] <= 32'b00001111000001100001000000000001;
REG[4061] <= 32'b11111100111110010000011011111010;
REG[4062] <= 32'b11111111111011011111000100000010;
REG[4063] <= 32'b11111101000100011111101111101101;
REG[4064] <= 32'b11110001111111001110111100001110;
REG[4065] <= 32'b00000000111101111110111100000110;
REG[4066] <= 32'b11111111000011000000000011110110;
REG[4067] <= 32'b11100111111100111111000000000001;
REG[4068] <= 32'b00001001111110111111011111110100;
REG[4069] <= 32'b11110001111110000000010111111010;
REG[4070] <= 32'b11110110111100011111010000000001;
REG[4071] <= 32'b11111101000000001111101000001000;
REG[4072] <= 32'b00001110000010101111101111111111;
REG[4073] <= 32'b11111100000010000000100100010100;
REG[4074] <= 32'b11111111111111011111101111111101;
REG[4075] <= 32'b00001000000011000000010000001001;
REG[4076] <= 32'b00001001111101011111000011101111;
REG[4077] <= 32'b00001001000100110001100100000110;
REG[4078] <= 32'b11111010111110110000110100001110;
REG[4079] <= 32'b00100000000000011111001011111010;
REG[4080] <= 32'b11110100111111001111100100000101;
REG[4081] <= 32'b00011001000100011111101011111110;
REG[4082] <= 32'b11110111000000010011000100010110;
REG[4083] <= 32'b11111101111110101111100100000010;
REG[4084] <= 32'b00001111111101101111001111111100;
REG[4085] <= 32'b00000010111100000000010011110111;
REG[4086] <= 32'b00000000000010100001001011111110;
REG[4087] <= 32'b00001110111011111111000111110110;
REG[4088] <= 32'b11111101111111010000010111110101;
REG[4089] <= 32'b11111110000001010000001011111011;
REG[4090] <= 32'b11110100111110100000101000011101;
REG[4091] <= 32'b00100011000100101111110100000010;
REG[4092] <= 32'b11111001111001111111100000000100;
REG[4093] <= 32'b11111010111111001111110111101010;
REG[4094] <= 32'b00000101111110110000000011110111;
REG[4095] <= 32'b11110011110111011110001100001110;
REG[4096] <= 32'b11110110000001011111100011110011;
REG[4097] <= 32'b00000000000010101111111000000111;
REG[4098] <= 32'b11110110111011011111110000000010;
REG[4099] <= 32'b00001000111110010000100000010010;
REG[4100] <= 32'b00000000111111100001001000000110;
REG[4101] <= 32'b11111100111101100000100111110110;
REG[4102] <= 32'b00001001111100100000011111110110;
REG[4103] <= 32'b00000001000001101111001100000101;
REG[4104] <= 32'b11110100111011011111111111111010;
REG[4105] <= 32'b11101111000100101110111111110100;
REG[4106] <= 32'b00001011111101111111001100001010;
REG[4107] <= 32'b11110101111101100000010011110000;
REG[4108] <= 32'b11101010111101011111011000000001;
REG[4109] <= 32'b00001011111101101111001111101001;
REG[4110] <= 32'b11110010111110010000001100000000;
REG[4111] <= 32'b11111001111101111111001111110000;
REG[4112] <= 32'b11110000111101101111100011110100;
REG[4113] <= 32'b11101100111100001111100011111010;
REG[4114] <= 32'b11110111111110101111101111111001;
REG[4115] <= 32'b11101101111110001111011111110100;
REG[4116] <= 32'b11111100111110001111010011111110;
REG[4117] <= 32'b11110111000001000000000011110101;
REG[4118] <= 32'b11110111000000101111100100000011;
REG[4119] <= 32'b00000010111101011111110100000000;
REG[4120] <= 32'b11111111000000110000100000000010;
REG[4121] <= 32'b11111110111111010000011111100101;
REG[4122] <= 32'b00001010000000110000100100000111;
REG[4123] <= 32'b01001100111001001111110111111110;
REG[4124] <= 32'b00010100111100100000001011100000;
REG[4125] <= 32'b00000010111100111111001011110000;
REG[4126] <= 32'b11111010111110010000011011110111;
REG[4127] <= 32'b11111000000101000001111011111011;
REG[4128] <= 32'b00000110000001000000001000001010;
REG[4129] <= 32'b00001111000001000001000100001000;
REG[4130] <= 32'b11111000000000011111110100000010;
REG[4131] <= 32'b00001000000011100000101100000111;
REG[4132] <= 32'b00000000111101000000001111111011;
REG[4133] <= 32'b11111111000000000000110111111011;
REG[4134] <= 32'b11111001111111100000011000000011;
REG[4135] <= 32'b11101000111010110000000011111100;
REG[4136] <= 32'b11111011000001011110011111100110;
REG[4137] <= 32'b00000110000011100000111000001010;
REG[4138] <= 32'b11101111111100011111001111111111;
REG[4139] <= 32'b00000110111111101110111111111001;
REG[4140] <= 32'b11111101000011010000100000000000;
REG[4141] <= 32'b11110110111011011111011100001011;
REG[4142] <= 32'b00000011111110101111111011110111;
REG[4143] <= 32'b00001000000000000000001011101000;
REG[4144] <= 32'b11110110111011000000010000000000;
REG[4145] <= 32'b00000011111011111111011111111011;
REG[4146] <= 32'b00000001111110111111111011101010;
REG[4147] <= 32'b11101110111101001111100011110010;
REG[4148] <= 32'b11110000111111001110111011101100;
REG[4149] <= 32'b11110001111110011111001000000110;
REG[4150] <= 32'b11111111111111101111001011110001;
REG[4151] <= 32'b11110000000001101111101111111110;
REG[4152] <= 32'b11111000000001000001000011110100;
REG[4153] <= 32'b00000110111100001111110011111101;
REG[4154] <= 32'b11111101000011000100100000010100;
REG[4155] <= 32'b00000000000001110000101111110111;
REG[4156] <= 32'b00001000111111010000011011111101;
REG[4157] <= 32'b11110110000010000000100000000011;
REG[4158] <= 32'b00000101000001000001000111111101;
REG[4159] <= 32'b11111100000000011111111111110011;
REG[4160] <= 32'b11111110000010111111101111110101;
REG[4161] <= 32'b11101111000101100001100111110100;
REG[4162] <= 32'b11101110111101111111010000101100;
REG[4163] <= 32'b00111100111010001110110000000001;
REG[4164] <= 32'b11110011000011010000100011110111;
REG[4165] <= 32'b11110110000001110000011100001000;
REG[4166] <= 32'b11111111000000110000100100000000;
REG[4167] <= 32'b00001010000000111111110100010000;
REG[4168] <= 32'b00000001111011111111101011110111;
REG[4169] <= 32'b00000010000000010000010111101010;
REG[4170] <= 32'b00001100000001001111101011111010;
REG[4171] <= 32'b11110001000000110000000011101000;
REG[4172] <= 32'b11101110111101011111001011111011;
REG[4173] <= 32'b11101001111000101110100111111010;
REG[4174] <= 32'b11110111111110001111100111111101;
REG[4175] <= 32'b11101111111111111111111000001001;
REG[4176] <= 32'b00101000001001110001101011110110;
REG[4177] <= 32'b11110010111111011111111111101001;
REG[4178] <= 32'b11110111111111111111111011111010;
REG[4179] <= 32'b11111111000000100000011000000000;
REG[4180] <= 32'b00001111000001010000001000000001;
REG[4181] <= 32'b00000011000010010001101100001010;
REG[4182] <= 32'b00000001111111011111111100010110;
REG[4183] <= 32'b00100111000101010000100100001110;
REG[4184] <= 32'b00001101000000011111101100000000;
REG[4185] <= 32'b11111111000100110000110111111001;
REG[4186] <= 32'b11110100111111101111010000000010;
REG[4187] <= 32'b00000000111110011110110111110110;
REG[4188] <= 32'b00001110111111111111010111101011;
REG[4189] <= 32'b11110101111100100000010100001010;
REG[4190] <= 32'b00000000111100101111000111110011;
REG[4191] <= 32'b00001100000000100000100011110000;
REG[4192] <= 32'b11110001111011000000000000001110;
REG[4193] <= 32'b00101010000001110000010000001010;
REG[4194] <= 32'b11111001111100100000111000000110;
REG[4195] <= 32'b11111100111111010000000111110100;
REG[4196] <= 32'b11110100111101100000110100000101;
REG[4197] <= 32'b00000111000000011111101111111100;
REG[4198] <= 32'b11110111111100110001010000000010;
REG[4199] <= 32'b11111100111011011111010111110100;
REG[4200] <= 32'b00010111000001100000011111111000;
REG[4201] <= 32'b11110011111101110000110011101100;
REG[4202] <= 32'b11110001111110100000010000010011;
REG[4203] <= 32'b00010001000010011110110011111100;
REG[4204] <= 32'b11110101000011001111110011110001;
REG[4205] <= 32'b11100110000000011111011000001110;
REG[4206] <= 32'b11111111000010100001001111101111;
REG[4207] <= 32'b11110000111101011111111100001000;
REG[4208] <= 32'b00000010111111011111011111111000;
REG[4209] <= 32'b00000000000000101110100111110011;
REG[4210] <= 32'b11101001111011011111011011111000;
REG[4211] <= 32'b11111101111111001111100100001011;
REG[4212] <= 32'b11101011000000011111011111111111;
REG[4213] <= 32'b00001000000101001111000000010101;
REG[4214] <= 32'b11111010111111000000100000010001;
REG[4215] <= 32'b11110110111110011111101011101101;
REG[4216] <= 32'b11101101111011000000001111110000;
REG[4217] <= 32'b11110101111011001111000111110010;
REG[4218] <= 32'b00001010111111001111101111101010;
REG[4219] <= 32'b11110000111011101111100111111011;
REG[4220] <= 32'b11111000000011101111100011111110;
REG[4221] <= 32'b11111100111101101111101100001100;
REG[4222] <= 32'b11111101000001011111101111101110;
REG[4223] <= 32'b11110111000011001111111111111110;
REG[4224] <= 32'b11111010000000011111101011111001;
REG[4225] <= 32'b00000110000010101111100011111000;
REG[4226] <= 32'b11110110111101000000010000001010;
REG[4227] <= 32'b11111011111110010000000011111101;
REG[4228] <= 32'b11111110000010111111000111101110;
REG[4229] <= 32'b11101011111110000000001111111100;
REG[4230] <= 32'b11110010111101011110111011111001;
REG[4231] <= 32'b11111011111101101111100111110100;
REG[4232] <= 32'b11110010111101101111010011111100;
REG[4233] <= 32'b00001101000001001111110011101100;
REG[4234] <= 32'b11110111111111100010010000001011;
REG[4235] <= 32'b00000001111100111111011011111101;
REG[4236] <= 32'b00000011111110111110011111110101;
REG[4237] <= 32'b11111000000001010000000100000101;
REG[4238] <= 32'b11111101000001101110101011101101;
REG[4239] <= 32'b11111110111111111111010000011111;
REG[4240] <= 32'b00100101000100101111110100000011;
REG[4241] <= 32'b00000001111110111111110100000110;
REG[4242] <= 32'b11110101111111110000001011111100;
REG[4243] <= 32'b11111010000000010001000100010111;
REG[4244] <= 32'b00010000000010000000001111111001;
REG[4245] <= 32'b00001001000011010000100100001010;
REG[4246] <= 32'b00000001111111100000111100010000;
REG[4247] <= 32'b00001100111101001111010011111100;
REG[4248] <= 32'b00000001111111000000110111111001;
REG[4249] <= 32'b00000001000011100000100000000011;
REG[4250] <= 32'b00000101111111100000001000010110;
REG[4251] <= 32'b11110101000000101111110111111001;
REG[4252] <= 32'b00000100000001011111110111111111;
REG[4253] <= 32'b11111001111110000000100000010001;
REG[4254] <= 32'b11111011111111100000001011111000;
REG[4255] <= 32'b00000111000010111111110000001001;
REG[4256] <= 32'b00000100111011101111100111101010;
REG[4257] <= 32'b00001011000100000001010111111110;
REG[4258] <= 32'b11111101111010010000001100000101;
REG[4259] <= 32'b00001010111111011111111111110010;
REG[4260] <= 32'b11110010111011101111110111111011;
REG[4261] <= 32'b11100110000000101110110011110010;
REG[4262] <= 32'b00000000111001111101100000000001;
REG[4263] <= 32'b11111100111101010000011100010000;
REG[4264] <= 32'b00000011000011100000001011110000;
REG[4265] <= 32'b00001001111101100000000000000011;
REG[4266] <= 32'b00000000111100110000101000000001;
REG[4267] <= 32'b11110111111111110000000000001110;
REG[4268] <= 32'b11111001111110100000011000001010;
REG[4269] <= 32'b11111011111111001111010011111100;
REG[4270] <= 32'b11111011111110101111100111111011;
REG[4271] <= 32'b11111001000001100000100011111001;
REG[4272] <= 32'b11110011111110110000011000001011;
REG[4273] <= 32'b00000110111110011111011011111000;
REG[4274] <= 32'b00000100111110010000100100000111;
REG[4275] <= 32'b11111101111110110000011100000001;
REG[4276] <= 32'b00010110000011011111110100000100;
REG[4277] <= 32'b00000111000001110000111000000010;
REG[4278] <= 32'b00000010111110101111111111111100;
REG[4279] <= 32'b11111110000000010000010100000111;
REG[4280] <= 32'b11111111111100011111000111110111;
REG[4281] <= 32'b11110011111110110000001000000001;
REG[4282] <= 32'b11110111111101110000010000000011;
REG[4283] <= 32'b11111100111110111111101000000010;
REG[4284] <= 32'b11110011111110111111100100000110;
REG[4285] <= 32'b11111001111111010000001100001001;
REG[4286] <= 32'b11111110000010101111101000000111;
REG[4287] <= 32'b00001011000001111111011100001010;
REG[4288] <= 32'b00001011000000000000101111111110;
REG[4289] <= 32'b11110011000111100010000000001011;
REG[4290] <= 32'b00010001000000011111100000010001;
REG[4291] <= 32'b00000111111110110000011100001011;
REG[4292] <= 32'b00000011111111111111101100000100;
REG[4293] <= 32'b00000101000101010000010000001001;
REG[4294] <= 32'b11111101111110000000011100000110;
REG[4295] <= 32'b11110111111110101111101011110011;
REG[4296] <= 32'b11111001111111000000100111111110;
REG[4297] <= 32'b11111011111101001111000011111110;
REG[4298] <= 32'b00000111111111100000100011101101;
REG[4299] <= 32'b11110111000001010000111100000001;
REG[4300] <= 32'b00001011111111101111101111111111;
REG[4301] <= 32'b00000111111110000000010111111011;
REG[4302] <= 32'b11110011111011110000010111110100;
REG[4303] <= 32'b00010001000011001111101111110011;
REG[4304] <= 32'b11111000000001100001001100010000;
REG[4305] <= 32'b00000000000100101111001111110111;
REG[4306] <= 32'b11110011000001010000011100010110;
REG[4307] <= 32'b11110111000001011111010100000001;
REG[4308] <= 32'b00000111000011101111100100000010;
REG[4309] <= 32'b11101110000000101111010011110100;
REG[4310] <= 32'b11111010111110001111000011111111;
REG[4311] <= 32'b11101110111100011110111111111000;
REG[4312] <= 32'b11110011000011100000011011111100;
REG[4313] <= 32'b00000011000000011111101100001010;
REG[4314] <= 32'b11110100111011111111001000000100;
REG[4315] <= 32'b11111111000001011111001111110000;
REG[4316] <= 32'b11110100111110111111100111111010;
REG[4317] <= 32'b11111010111110001111101011110011;
REG[4318] <= 32'b11110100111110100000001111111111;
REG[4319] <= 32'b11111010111111000000100100000111;
REG[4320] <= 32'b11110111111101001111110111111010;
REG[4321] <= 32'b11111111000000010000010100000010;
REG[4322] <= 32'b11111101111101111110110011110010;
REG[4323] <= 32'b00000000000000001111100100000111;
REG[4324] <= 32'b11111110111101010000101111111111;
REG[4325] <= 32'b11111100000001011111111011110100;
REG[4326] <= 32'b11110111111100111111101100000111;
REG[4327] <= 32'b00001000000000101111010111110110;
REG[4328] <= 32'b11111000000010011111100111101110;
REG[4329] <= 32'b11111001111101001111100100010001;
REG[4330] <= 32'b00000110000101101111011111111010;
REG[4331] <= 32'b11111000000011010000011100010010;
REG[4332] <= 32'b00000100111101001111001100000111;
REG[4333] <= 32'b11111110111110100000010111111110;
REG[4334] <= 32'b11111111111101001111111111110110;
REG[4335] <= 32'b00000001111110010000011111110001;
REG[4336] <= 32'b11110111111011101111011011011111;
REG[4337] <= 32'b11110101000011110000010011111101;
REG[4338] <= 32'b11110110110111111110100000010111;
REG[4339] <= 32'b00001011111110100000100011101010;
REG[4340] <= 32'b11110110111111100000000100000000;
REG[4341] <= 32'b00000001000010010000000100000011;
REG[4342] <= 32'b11111100000010100000011000010001;
REG[4343] <= 32'b00001110111111101111110100000110;
REG[4344] <= 32'b00000101000010100001000011111100;
REG[4345] <= 32'b11111000111111011111110011111101;
REG[4346] <= 32'b00010011000011110000100100000001;
REG[4347] <= 32'b11111000111110001111101111111000;
REG[4348] <= 32'b00000001111110110000000100000000;
REG[4349] <= 32'b00000100000001100001010100001100;
REG[4350] <= 32'b00010010000000011111000011111010;
REG[4351] <= 32'b00000101111111010000011111111000;
REG[4352] <= 32'b00000000111101110001100011111101;
REG[4353] <= 32'b11111110111100001111000111111110;
REG[4354] <= 32'b00001110111111000000101100000001;
REG[4355] <= 32'b00001011000000001111110011110111;
REG[4356] <= 32'b11111011111101000000000011110111;
REG[4357] <= 32'b11111011000000111111111100000000;
REG[4358] <= 32'b11111100111100000000001000011110;
REG[4359] <= 32'b00010111000010001111100011111011;
REG[4360] <= 32'b00100010000000000010011000010000;
REG[4361] <= 32'b11110111111110010010010011110110;
REG[4362] <= 32'b00101000000101111111111011110011;
REG[4363] <= 32'b00100001111110101111100011110100;
REG[4364] <= 32'b00000000111011111111001111111001;
REG[4365] <= 32'b11111010111101001111101111110010;
REG[4366] <= 32'b11110101111111111111111011111011;
REG[4367] <= 32'b11111110111100101111011111111110;
REG[4368] <= 32'b11110101111110001111010011110011;
REG[4369] <= 32'b11110111000000011111000011111011;
REG[4370] <= 32'b11111100111101100000000100000010;
REG[4371] <= 32'b11101111111101011111001011111110;
REG[4372] <= 32'b00000101000000001110101011110011;
REG[4373] <= 32'b00010011111110101111111000000000;
REG[4374] <= 32'b11110101000110110010011111110110;
REG[4375] <= 32'b11111110111111001111000100011011;
REG[4376] <= 32'b00001101111101100000001011111010;
REG[4377] <= 32'b11111010111111110000001111111111;
REG[4378] <= 32'b11111100111110011111000011111010;
REG[4379] <= 32'b11111110000001011111100000001010;
REG[4380] <= 32'b11111011111110110000001111111101;
REG[4381] <= 32'b11110100111101010000110111111010;
REG[4382] <= 32'b00000111000011110000101000000000;
REG[4383] <= 32'b11111101111010000000100100001011;
REG[4384] <= 32'b11111101111101100000010011110110;
REG[4385] <= 32'b00001011111110110000000100000011;
REG[4386] <= 32'b11111111000001110000011011110011;
REG[4387] <= 32'b11111000111111010010000000001100;
REG[4388] <= 32'b00010011111011111111101011111110;
REG[4389] <= 32'b11101011111110011111100111110000;
REG[4390] <= 32'b11111010111111010000011000010010;
REG[4391] <= 32'b00010000000000111111110000001010;
REG[4392] <= 32'b00000100000001111111111000001001;
REG[4393] <= 32'b00001010000011000000010111111110;
REG[4394] <= 32'b11111010111110011111101111111100;
REG[4395] <= 32'b11110110111101101111011000001000;
REG[4396] <= 32'b00111110001010001111011111111000;
REG[4397] <= 32'b00000111000011100100001000011011;
REG[4398] <= 32'b11111001111110110000010111111111;
REG[4399] <= 32'b00101000000000011111011111111101;
REG[4400] <= 32'b00010101000000000000000011111001;
REG[4401] <= 32'b11111001111111110001111100000100;
REG[4402] <= 32'b00000000111110011111001111110000;
REG[4403] <= 32'b00000001000001010000010000010001;
REG[4404] <= 32'b11111111111110110000010011100100;
REG[4405] <= 32'b11101110000001110000011100000010;
REG[4406] <= 32'b00000111111000111110110100000000;
REG[4407] <= 32'b00000000111111110000010011111000;
REG[4408] <= 32'b11110110111111001111011100001000;
REG[4409] <= 32'b11101101111111100000011100001101;
REG[4410] <= 32'b00010110000111011111100000010010;
REG[4411] <= 32'b11111111000000111111101111110011;
REG[4412] <= 32'b11101100000010100000010100000111;
REG[4413] <= 32'b11111101000001001111111011101000;
REG[4414] <= 32'b11101000111001011111111011111101;
REG[4415] <= 32'b11110110111101111110111111110001;
REG[4416] <= 32'b11111100111110001110111111111010;
REG[4417] <= 32'b11110001111011011110101011101011;
REG[4418] <= 32'b11101111111111011111100000000001;
REG[4419] <= 32'b11110110111111111111111000001011;
REG[4420] <= 32'b00001011111111111110111011110010;
REG[4421] <= 32'b11110010000000110000010100010000;
REG[4422] <= 32'b11111010000000100000000011111110;
REG[4423] <= 32'b11111101000000011111111011110010;
REG[4424] <= 32'b11110110000010100000011000000011;
REG[4425] <= 32'b00000011111111011111001011110110;
REG[4426] <= 32'b11111011111111000000010000000011;
REG[4427] <= 32'b00000010111111000000101100000101;
REG[4428] <= 32'b11110110111111101111101011110110;
REG[4429] <= 32'b00010000000001101111110011111011;
REG[4430] <= 32'b11111000000000100000111100000110;
REG[4431] <= 32'b00000110111101100000110111110111;
REG[4432] <= 32'b00001001000010100000001100000000;
REG[4433] <= 32'b00001101000010100001011000001010;
REG[4434] <= 32'b00011111000110010010110100001000;
REG[4435] <= 32'b00000110000010110000010100000110;
REG[4436] <= 32'b11111100000001010000010000000010;
REG[4437] <= 32'b11111001111110011111100011111011;
REG[4438] <= 32'b11111111111111011111001011110001;
REG[4439] <= 32'b11110111111111111111010111111110;
REG[4440] <= 32'b11110110111100001110111011101011;
REG[4441] <= 32'b11100100111001101111001111110100;
REG[4442] <= 32'b11101110111010001110010011100111;
REG[4443] <= 32'b11110010111101111111100111110110;
REG[4444] <= 32'b11101011111101000000010111111101;
REG[4445] <= 32'b00100000111101010000001000000001;
REG[4446] <= 32'b00001100000000010001100011110010;
REG[4447] <= 32'b00001111000100110001000100000010;
REG[4448] <= 32'b00001111111111101111110011110110;
REG[4449] <= 32'b11110010000000000000010111101111;
REG[4450] <= 32'b11111101000001111110100111111010;
REG[4451] <= 32'b00000001111100101111101011111110;
REG[4452] <= 32'b11111011000001010000010011110001;
REG[4453] <= 32'b11110110111110100000101100000000;
REG[4454] <= 32'b00000000000001010000010100001100;
REG[4455] <= 32'b00010101000001001111110000000000;
REG[4456] <= 32'b11111000111111000000101100000010;
REG[4457] <= 32'b00000000111101101111101011111010;
REG[4458] <= 32'b11110110111101001110100111111001;
REG[4459] <= 32'b11111001111101000000001111111101;
REG[4460] <= 32'b11110111111100101110111011101011;
REG[4461] <= 32'b11110001111110101111110011111100;
REG[4462] <= 32'b11111111111101110000000100000011;
REG[4463] <= 32'b00001111111101010000111000000101;
REG[4464] <= 32'b11111011111100110000101000001001;
REG[4465] <= 32'b00100100000111000000101000000110;
REG[4466] <= 32'b00001011000011010000010000000111;
REG[4467] <= 32'b00001111111110001111100111101111;
REG[4468] <= 32'b11101100111010010011000100000110;
REG[4469] <= 32'b00001001111001111110101111101101;
REG[4470] <= 32'b00001011111111001111110011100011;
REG[4471] <= 32'b11101010111100000000011000000100;
REG[4472] <= 32'b11110011000001011111011011111001;
REG[4473] <= 32'b00000110000000111111111000001010;
REG[4474] <= 32'b00000100000010010000000100000001;
REG[4475] <= 32'b11111011000010110000000011111010;
REG[4476] <= 32'b00001110000010101111111011101110;
REG[4477] <= 32'b11111011000001110000101000001100;
REG[4478] <= 32'b00000100111011111111100100000010;
REG[4479] <= 32'b00001110000011100000111011110011;
REG[4480] <= 32'b11111011111111111111011011111011;
REG[4481] <= 32'b00000001000011001111100111111110;
REG[4482] <= 32'b11110010111110010000001100000010;
REG[4483] <= 32'b11101011111100011111110011111001;
REG[4484] <= 32'b00000100000101100000011100000011;
REG[4485] <= 32'b11111100000000011111011111111101;
REG[4486] <= 32'b11111100111110000000011111111111;
REG[4487] <= 32'b11111101111110001111101011111000;
REG[4488] <= 32'b11110101000001000000000000000000;
REG[4489] <= 32'b11111101111101111111110111111101;
REG[4490] <= 32'b11111001000101100000011011110010;
REG[4491] <= 32'b11111011111110111111011100010001;
REG[4492] <= 32'b00000000111011011111100111111000;
REG[4493] <= 32'b11101010000100100000000111110101;
REG[4494] <= 32'b00000000000001000000001100000100;
REG[4495] <= 32'b00000010111110011111100000010010;
REG[4496] <= 32'b00000010111111101111111011111000;
REG[4497] <= 32'b11110110000011110000011000000101;
REG[4498] <= 32'b00000011111110111111101100000010;
REG[4499] <= 32'b11111111000000001111110100000111;
REG[4500] <= 32'b11111111000001011111100000001110;
REG[4501] <= 32'b00000101000010011111011000000010;
REG[4502] <= 32'b11110010111111111111011000000000;
REG[4503] <= 32'b00010001001010110001011011110111;
REG[4504] <= 32'b11101110111101011111101000001100;
REG[4505] <= 32'b11111001111110101111000111111000;
REG[4506] <= 32'b00010010000111000000110011111100;
REG[4507] <= 32'b11101010111110000000011100000110;
REG[4508] <= 32'b00000010111110111111101100000001;
REG[4509] <= 32'b00000111111111111111011011111111;
REG[4510] <= 32'b00001000111110100001000011111111;
REG[4511] <= 32'b11110111000001100000000111110101;
REG[4512] <= 32'b00000101000001000000000000000001;
REG[4513] <= 32'b11111100111011110000100100000000;
REG[4514] <= 32'b00000001000010000000000000000110;
REG[4515] <= 32'b00001011000000011111100100001011;
REG[4516] <= 32'b00001010001000010000010000010001;
REG[4517] <= 32'b11111100000001110000100100000011;
REG[4518] <= 32'b00010000000010101111101100100000;
REG[4519] <= 32'b00010101000110100000000011110101;
REG[4520] <= 32'b11111011000110100001011000001100;
REG[4521] <= 32'b11111111000011110000110011110000;
REG[4522] <= 32'b11110001111110100000010011111000;
REG[4523] <= 32'b00000000111111101111011000000000;
REG[4524] <= 32'b00000010111111100000100000000000;
REG[4525] <= 32'b11101100111101010000000011100100;
REG[4526] <= 32'b00001001111111000000010100001011;
REG[4527] <= 32'b11101010111000001111001011111111;
REG[4528] <= 32'b11110011000000000000011100000101;
REG[4529] <= 32'b00001010000001001111101000001111;
REG[4530] <= 32'b00001011000000001111001011111001;
REG[4531] <= 32'b00001101000000110000110100010000;
REG[4532] <= 32'b00000100111100001111111111111101;
REG[4533] <= 32'b00010000000011101111100111110101;
REG[4534] <= 32'b00000011111001111111001100000010;
REG[4535] <= 32'b00000011111011101111101000000000;
REG[4536] <= 32'b11111110111111001111110111110001;
REG[4537] <= 32'b11111011000000010000100111111110;
REG[4538] <= 32'b00001110111111000001000011111111;
REG[4539] <= 32'b11110101111111000000011111110101;
REG[4540] <= 32'b11111010111011100000000011111101;
REG[4541] <= 32'b11111101111101101111011111110010;
REG[4542] <= 32'b00001010000001010000000111110111;
REG[4543] <= 32'b11111001111110100000010011110101;
REG[4544] <= 32'b11110110000100010000101100001011;
REG[4545] <= 32'b11111111000000010000000000011100;
REG[4546] <= 32'b00010000111111100000001111111110;
REG[4547] <= 32'b00000011000110010001011100000101;
REG[4548] <= 32'b00000100000000101111100000000110;
REG[4549] <= 32'b00000000111101011111100011110101;
REG[4550] <= 32'b11111001111110011111010011111011;
REG[4551] <= 32'b00000101000000111111111111111110;
REG[4552] <= 32'b00001010001010000010011011111010;
REG[4553] <= 32'b00000111111101111111011011111100;
REG[4554] <= 32'b00010110000001111111011100000001;
REG[4555] <= 32'b11111000111110011111110000000100;
REG[4556] <= 32'b11111111000011110000110000000101;
REG[4557] <= 32'b11111101000010000000101111111100;
REG[4558] <= 32'b00000000111101011111010011111011;
REG[4559] <= 32'b00000001111111101111011111110101;
REG[4560] <= 32'b11110011111101101111110011101010;
REG[4561] <= 32'b11101000111010110000000011111010;
REG[4562] <= 32'b00001101111111011111101000000000;
REG[4563] <= 32'b00000100000000100000010111111011;
REG[4564] <= 32'b00001001000001110000001011111000;
REG[4565] <= 32'b11111110000010110001010000000011;
REG[4566] <= 32'b00000000111110101111101000000010;
REG[4567] <= 32'b00010111000010100000011011111000;
REG[4568] <= 32'b11110101000001110001111100001000;
REG[4569] <= 32'b11111010000000001111101100000011;
REG[4570] <= 32'b11110100111110100000001100010000;
REG[4571] <= 32'b00000100111110111110111100001011;
REG[4572] <= 32'b11111101000011101111110000001000;
REG[4573] <= 32'b11111111000011101111010011111011;
REG[4574] <= 32'b11111010000010101111110100001001;
REG[4575] <= 32'b11111010000010100000001011110011;
REG[4576] <= 32'b11111101111101101111110111111111;
REG[4577] <= 32'b00000000111110011111010111111001;
REG[4578] <= 32'b11110000111101111111101111111001;
REG[4579] <= 32'b11111000111100011111010011111110;
REG[4580] <= 32'b00000010111101001111001111111010;
REG[4581] <= 32'b00000000111101111111101111101000;
REG[4582] <= 32'b11110101111110011111110011111110;
REG[4583] <= 32'b00001111111001011110111111101011;
REG[4584] <= 32'b00001000111111110000101111110100;
REG[4585] <= 32'b00100001000001110001001100000000;
REG[4586] <= 32'b00000100000100010001100011111111;
REG[4587] <= 32'b00010010111111111111110100001001;
REG[4588] <= 32'b00000100000001011111001011111011;
REG[4589] <= 32'b11111010111110101111101111101010;
REG[4590] <= 32'b11110100111111010000010100000100;
REG[4591] <= 32'b00001101111100101111100011111001;
REG[4592] <= 32'b00000001111111000000101111110011;
REG[4593] <= 32'b11101110111110100000001000001101;
REG[4594] <= 32'b00010100000001001111100000000001;
REG[4595] <= 32'b11111101000101000001011011111101;
REG[4596] <= 32'b11110111000001100000011100100001;
REG[4597] <= 32'b00100110111111000000110000000111;
REG[4598] <= 32'b11111100111110101111010111110111;
REG[4599] <= 32'b11110010000001111111111111111110;
REG[4600] <= 32'b11110111111110001111001100001100;
REG[4601] <= 32'b00000100000001110000001111111001;
REG[4602] <= 32'b11111110000001000000010100001100;
REG[4603] <= 32'b00001010000011101111011111111000;
REG[4604] <= 32'b11111001000010110000010100000101;
REG[4605] <= 32'b11111111111110111111101011111011;
REG[4606] <= 32'b11111100111110111111011100011100;
REG[4607] <= 32'b00100001000100110000010011110100;
REG[4608] <= 32'b00011101000101000000100100001011;
REG[4609] <= 32'b11111101111100111110110111101101;
REG[4610] <= 32'b11111000000001011111111111110001;
REG[4611] <= 32'b00000000000011010000000000001101;
REG[4612] <= 32'b00001000000001100000001000000100;
REG[4613] <= 32'b00000001000100000001011100000111;
REG[4614] <= 32'b00000110000011010000110100001110;
REG[4615] <= 32'b00010110000011000000000100001000;
REG[4616] <= 32'b11111011111101100000000100001000;
REG[4617] <= 32'b00001001000011000000000011111000;
REG[4618] <= 32'b00000001111110010000111011111111;
REG[4619] <= 32'b00000111111111000000011011111000;
REG[4620] <= 32'b00000001000000110000001111111111;
REG[4621] <= 32'b11111100111101110001001100011111;
REG[4622] <= 32'b00001011111101111111011111111000;
REG[4623] <= 32'b00001010000011110000101111111011;
REG[4624] <= 32'b11111010111110111111100000000001;
REG[4625] <= 32'b00001101111101010000001000001110;
REG[4626] <= 32'b11111001000101000001000111111101;
REG[4627] <= 32'b11111111111110110010101100011111;
REG[4628] <= 32'b11110001111100101111010011110011;
REG[4629] <= 32'b11111100111111010000110100011000;
REG[4630] <= 32'b11110011111010010000000111111101;
REG[4631] <= 32'b00001001000101000001000011101110;
REG[4632] <= 32'b00000010000000100000100011111010;
REG[4633] <= 32'b11110100111100010000000000001111;
REG[4634] <= 32'b00001001111110110000101100000100;
REG[4635] <= 32'b00001011000001001111100100000011;
REG[4636] <= 32'b00000011111110110000011000000000;
REG[4637] <= 32'b11110110000100111111100011110000;
REG[4638] <= 32'b11110000000001000010000100001110;
REG[4639] <= 32'b00001000111100011110111111110100;
REG[4640] <= 32'b11111010000010010000011011110111;
REG[4641] <= 32'b11111010111101101111101111110111;
REG[4642] <= 32'b11111101111011100000001000001000;
REG[4643] <= 32'b00001100000000111111100100001100;
REG[4644] <= 32'b11110100000010100000101100001001;
REG[4645] <= 32'b00001100000100001111111100001100;
REG[4646] <= 32'b11111100000010100001100100010001;
REG[4647] <= 32'b00001011000010001111011000001101;
REG[4648] <= 32'b00010001000100000000100100001110;
REG[4649] <= 32'b11110111000000100000100100000110;
REG[4650] <= 32'b00000010111111011111000100001001;
REG[4651] <= 32'b00000010111111111111101011110110;
REG[4652] <= 32'b11111000111111010000101000001110;
REG[4653] <= 32'b00000101111110101111101011101110;
REG[4654] <= 32'b00001000000100111111101011111111;
REG[4655] <= 32'b11111011111011010000100100010011;
REG[4656] <= 32'b00000110000000011111001011111000;
REG[4657] <= 32'b11101111000001010000000100000101;
REG[4658] <= 32'b11111101000000101111111000010110;
REG[4659] <= 32'b00000011000000001111100011111100;
REG[4660] <= 32'b11110111000000011111101011111110;
REG[4661] <= 32'b11111001111111110000101100000011;
REG[4662] <= 32'b11111110000000011111001000000010;
REG[4663] <= 32'b00000111000010011111101011111101;
REG[4664] <= 32'b11111010111111100000000100001110;
REG[4665] <= 32'b11111010000000101111010011110111;
REG[4666] <= 32'b11101111000101110000101011111111;
REG[4667] <= 32'b11111100000010011111000000001010;
REG[4668] <= 32'b11111000111111111111110111110010;
REG[4669] <= 32'b11110111000011011111101100000001;
REG[4670] <= 32'b00010110111011101111100000001000;
REG[4671] <= 32'b11110100111101010000000111110000;
REG[4672] <= 32'b11101001111100001111101100010100;
REG[4673] <= 32'b00100111111110011111011100000011;
REG[4674] <= 32'b00000110111100001111011111110101;
REG[4675] <= 32'b11110100111111110000000011110101;
REG[4676] <= 32'b11111100111101001111100011111100;
REG[4677] <= 32'b11110110111110010000100111110000;
REG[4678] <= 32'b11110110111101111111010111100111;
REG[4679] <= 32'b11101110111101101111010000000001;
REG[4680] <= 32'b11110110111101111110111011101111;
REG[4681] <= 32'b11101111111110001111010111101111;
REG[4682] <= 32'b11101101111110001111100011111101;
REG[4683] <= 32'b11110011000000000000010100001100;
REG[4684] <= 32'b00000000111111101111011011111000;
REG[4685] <= 32'b11111001000000001111011011110100;
REG[4686] <= 32'b00000111000001001111110111111110;
REG[4687] <= 32'b00000000111100111111100000000101;
REG[4688] <= 32'b11111101111110111111101111111000;
REG[4689] <= 32'b11110011111111101111100000001000;
REG[4690] <= 32'b00000000111110101110111111111001;
REG[4691] <= 32'b11110110000011010000011111110100;
REG[4692] <= 32'b00001100111111001111111000001100;
REG[4693] <= 32'b00000100000000101111010111101001;
REG[4694] <= 32'b11110010000001001111011000000100;
REG[4695] <= 32'b00000011111100011111110011111001;
REG[4696] <= 32'b11110001111111011111100011111110;
REG[4697] <= 32'b00001100111101101111010100011001;
REG[4698] <= 32'b11111001111111100000111011101000;
REG[4699] <= 32'b11111001111010001111111111111011;
REG[4700] <= 32'b11111100111101110000101100000100;
REG[4701] <= 32'b11111101111101011111100011111001;
REG[4702] <= 32'b11101001111011001111011011101001;
REG[4703] <= 32'b11101101111111100000111011111100;
REG[4704] <= 32'b00000100111100011111000000000010;
REG[4705] <= 32'b00101011000011011111110011111010;
REG[4706] <= 32'b00000000000001010000000011110101;
REG[4707] <= 32'b00000000111101100000001011101110;
REG[4708] <= 32'b11110111111110000000000111110010;
REG[4709] <= 32'b11110100000000000000000011101011;
REG[4710] <= 32'b11101111111100001111011011110100;
REG[4711] <= 32'b11111010000101011110111011101111;
REG[4712] <= 32'b11110101111111110000101100011011;
REG[4713] <= 32'b11110100111101101111010111101011;
REG[4714] <= 32'b11111001000001010000011100100100;
REG[4715] <= 32'b00010101000000111111010011110100;
REG[4716] <= 32'b00000011000101110000100100000110;
REG[4717] <= 32'b11111101000000001111100000000000;
REG[4718] <= 32'b11110010000001110000110100001011;
REG[4719] <= 32'b00001010000000110000000100000001;
REG[4720] <= 32'b11111100000001100000001100001100;
REG[4721] <= 32'b00001101111110001111001000000010;
REG[4722] <= 32'b00000011000011110000001011111001;
REG[4723] <= 32'b11101110000000100001101011111011;
REG[4724] <= 32'b00000000111011001110100011101110;
REG[4725] <= 32'b00001111111100001111000011110100;
REG[4726] <= 32'b11101010111011100001111111111100;
REG[4727] <= 32'b11111011000001100000000000000100;
REG[4728] <= 32'b11110000111101100000001111111011;
REG[4729] <= 32'b00001100000001110000011100100110;
REG[4730] <= 32'b00010011111101110000010000000010;
REG[4731] <= 32'b11111100000111110001101011111101;
REG[4732] <= 32'b00001011111101110000010011101011;
REG[4733] <= 32'b11110011000010100001101100010011;
REG[4734] <= 32'b00001000111100101110111011111011;
REG[4735] <= 32'b00001010111110111111101011100111;
REG[4736] <= 32'b11101001000000000000011111111110;
REG[4737] <= 32'b11110111111111110000101111111000;
REG[4738] <= 32'b11110010111110000000010000000001;
REG[4739] <= 32'b00001011111101001111001100000010;
REG[4740] <= 32'b11111110111101001111110111110100;
REG[4741] <= 32'b11110101000000010000001011111101;
REG[4742] <= 32'b11101101000010100000101100011001;
REG[4743] <= 32'b11111101111101011110010111110101;
REG[4744] <= 32'b11111110111110100000000111111001;
REG[4745] <= 32'b11101101111110111111111100000000;
REG[4746] <= 32'b00001000111111110000010100001001;
REG[4747] <= 32'b00101001111110000000001111111101;
REG[4748] <= 32'b00000010000001110001001100000010;
REG[4749] <= 32'b00000001000000110000001100010001;
REG[4750] <= 32'b11100101111011111111111111111001;
REG[4751] <= 32'b00000010001001000010000011011011;
REG[4752] <= 32'b11111100111110001111110100100010;
REG[4753] <= 32'b01010000111010000000000011111101;
REG[4754] <= 32'b00000001000010110001110000000000;
REG[4755] <= 32'b11111101000000100000011011111010;
REG[4756] <= 32'b11111101000000110000010100001011;
REG[4757] <= 32'b00000100111111000000100100001110;
REG[4758] <= 32'b00000110000001011111101011111101;
REG[4759] <= 32'b00010000000001100000011111111101;
REG[4760] <= 32'b00000100000001001111110000001010;
REG[4761] <= 32'b11110111111101000000101100001101;
REG[4762] <= 32'b11111001111110100000100100000100;
REG[4763] <= 32'b00010000000100011111110100000110;
REG[4764] <= 32'b11110001111101110000000011110100;
REG[4765] <= 32'b00000011111101111111101111111011;
REG[4766] <= 32'b11111001111100111111101011110100;
REG[4767] <= 32'b11111011111011111111110011101000;
REG[4768] <= 32'b11110110111110010001001000010010;
REG[4769] <= 32'b00000000000001001111000011110110;
REG[4770] <= 32'b00001100001110010001001000000111;
REG[4771] <= 32'b00010011111110010001000100001101;
REG[4772] <= 32'b00000010000101000001101100010000;
REG[4773] <= 32'b11111100000001010000011011110010;
REG[4774] <= 32'b11111100000101011111011000001111;
REG[4775] <= 32'b00000001111110110000000000001000;
REG[4776] <= 32'b00000100000101100000100000001101;
REG[4777] <= 32'b00010010000110100000100011111001;
REG[4778] <= 32'b00001111111110011111001111111101;
REG[4779] <= 32'b11111111111111000000110100001000;
REG[4780] <= 32'b00000111000100101111111111111100;
REG[4781] <= 32'b00010001000010000000001100000101;
REG[4782] <= 32'b11111101111101110000101011110110;
REG[4783] <= 32'b11111000111111010000001111111110;
REG[4784] <= 32'b11111100111100110000010000000100;
REG[4785] <= 32'b11111111111110001111000011110001;
REG[4786] <= 32'b11111111000000101111011111111010;
REG[4787] <= 32'b00000000000011110000111100000011;
REG[4788] <= 32'b11110011111101111111101011110001;
REG[4789] <= 32'b11110110111011111111010111111100;
REG[4790] <= 32'b11110110111110000000001000001000;
REG[4791] <= 32'b11111100111100101111011111111101;
REG[4792] <= 32'b11110101111110011111101111111001;
REG[4793] <= 32'b11111100111111101111100011111101;
REG[4794] <= 32'b11111010111100111111001000000111;
REG[4795] <= 32'b11110111000000001110010111100111;
REG[4796] <= 32'b11110110111101101111001111110010;
REG[4797] <= 32'b11100111111011101111010011111101;
REG[4798] <= 32'b11110001111101001110011111101011;
REG[4799] <= 32'b11110111000000111111101000000010;
REG[4800] <= 32'b11111101000000110000100000001001;
REG[4801] <= 32'b11111111000010100000010000001101;
REG[4802] <= 32'b11111010000011000000011000010100;
REG[4803] <= 32'b11110110111100111111000000000000;
REG[4804] <= 32'b00000011000010100000011011111011;
REG[4805] <= 32'b00001011000001000001000011111001;
REG[4806] <= 32'b00000000111101001111011100000101;
REG[4807] <= 32'b00000110111101101111011011111101;
REG[4808] <= 32'b11111010000001110000000011111110;
REG[4809] <= 32'b00001011111011111111010111111110;
REG[4810] <= 32'b11100010111100100000111011110011;
REG[4811] <= 32'b11110010111100111111110000000101;
REG[4812] <= 32'b00000011111100001111001000000011;
REG[4813] <= 32'b00010010000010111111110111111110;
REG[4814] <= 32'b00000011111100011111010000000010;
REG[4815] <= 32'b00001000111110111111101111111100;
REG[4816] <= 32'b00000011000011110000110011111011;
REG[4817] <= 32'b00000001111110101111110100001010;
REG[4818] <= 32'b11111010111100011111010100000001;
REG[4819] <= 32'b00000110111101111111110011110011;
REG[4820] <= 32'b00010010000001111111110111110110;
REG[4821] <= 32'b11110001111101100000110111111011;
REG[4822] <= 32'b11110101111011111111101111110111;
REG[4823] <= 32'b11111000000000111111111100000010;
REG[4824] <= 32'b11111100000000101111010100000110;
REG[4825] <= 32'b11111100000001001111010000000101;
REG[4826] <= 32'b00000101111011101111101011111110;
REG[4827] <= 32'b11110001000010000001010000001010;
REG[4828] <= 32'b00001011111101111111011100001001;
REG[4829] <= 32'b00010010111111101111101111101100;
REG[4830] <= 32'b11111100111110100000000111110001;
REG[4831] <= 32'b11110110111101001111100100000100;
REG[4832] <= 32'b00000101000001001111011011111101;
REG[4833] <= 32'b11110111111111111111110100000011;
REG[4834] <= 32'b00000001000000110000000100000001;
REG[4835] <= 32'b00000001111111011111100111110011;
REG[4836] <= 32'b00000010111101000000001111101111;
REG[4837] <= 32'b00000111000111100000100011111001;
REG[4838] <= 32'b11111100111100110000111000011001;
REG[4839] <= 32'b11110001111100001111111011110011;
REG[4840] <= 32'b00000011000000101111011011111101;
REG[4841] <= 32'b11101101111110101110101000000101;
REG[4842] <= 32'b00000110000111001111001000000011;
REG[4843] <= 32'b11101111000010001111110100001101;
REG[4844] <= 32'b11111000000101000000101000010100;
REG[4845] <= 32'b00000110000001011111110111110000;
REG[4846] <= 32'b11111000111111010001010000000000;
REG[4847] <= 32'b00000101000001001111010011110011;
REG[4848] <= 32'b00000001000000100001000000000111;
REG[4849] <= 32'b00000111000010011111111111111100;
REG[4850] <= 32'b00000010111111011111001011110110;
REG[4851] <= 32'b00001101111111011111111011111010;
REG[4852] <= 32'b11110011111101010000100100001001;
REG[4853] <= 32'b00000011111110101111010011111101;
REG[4854] <= 32'b11110101111110001111110000010100;
REG[4855] <= 32'b00001011111101101111010011111100;
REG[4856] <= 32'b11111011000100110000111011111100;
REG[4857] <= 32'b11111001000000011111010000000100;
REG[4858] <= 32'b11111011111010100000000111111011;
REG[4859] <= 32'b00000000111100111111110011101111;
REG[4860] <= 32'b11110111111101001111100111110010;
REG[4861] <= 32'b11111001111010101111110011111101;
REG[4862] <= 32'b11111000000000001111101011110110;
REG[4863] <= 32'b11110010111110001111110111110111;
REG[4864] <= 32'b11110111111011001111101011111000;
REG[4865] <= 32'b11110100111111101111111011110011;
REG[4866] <= 32'b11111000111110101111111011111111;
REG[4867] <= 32'b11111110111101110000000100000010;
REG[4868] <= 32'b00010000000000110000001000011111;
REG[4869] <= 32'b00000000000000101111110100000110;
REG[4870] <= 32'b00000000000110101111111100000010;
REG[4871] <= 32'b11111001000011000000110000001111;
REG[4872] <= 32'b00000111000000100000010100000000;
REG[4873] <= 32'b11111100111111101111001111100101;
REG[4874] <= 32'b11110011000111000001010011111101;
REG[4875] <= 32'b11111100111110001111111111111011;
REG[4876] <= 32'b11110010111101101111100100000000;
REG[4877] <= 32'b11110111000010101111101011110111;
REG[4878] <= 32'b00001001000000101111010000001011;
REG[4879] <= 32'b11110101111101100001100100010101;
REG[4880] <= 32'b11110001111111111111000111101101;
REG[4881] <= 32'b00001100000000001111010100011100;
REG[4882] <= 32'b00010001111110001111010000001000;
REG[4883] <= 32'b00000100000101010000011011111001;
REG[4884] <= 32'b11110010111110000000001000001110;
REG[4885] <= 32'b11101101111010101111000111101100;
REG[4886] <= 32'b11111010111011011111010111111010;
REG[4887] <= 32'b00001101111011111111100011110011;
REG[4888] <= 32'b11111001111110010010001000001011;
REG[4889] <= 32'b11110001111011011111101111111010;
REG[4890] <= 32'b11111101111110101111010100001100;
REG[4891] <= 32'b00001000111101011111010111110101;
REG[4892] <= 32'b11110110001000000010001000000011;
REG[4893] <= 32'b00001001111110101111110011011011;
REG[4894] <= 32'b11101111111001011111101000000000;
REG[4895] <= 32'b11110101000010110000010000001100;
REG[4896] <= 32'b11110111111111111111110100010001;
REG[4897] <= 32'b11111110111110011111110011111110;
REG[4898] <= 32'b11111000000010101111110011110010;
REG[4899] <= 32'b11110001111110100000000111111000;
REG[4900] <= 32'b00000011000001011111001111111010;
REG[4901] <= 32'b00000011111110101111011100000000;
REG[4902] <= 32'b00000001000000010000001111110101;
REG[4903] <= 32'b11110000111100111111010111111100;
REG[4904] <= 32'b00001110000001000000100100000010;
REG[4905] <= 32'b11110010111110100000101000000110;
REG[4906] <= 32'b11111100000010001111000011111000;
REG[4907] <= 32'b00000001111100111111001011101100;
REG[4908] <= 32'b11110010111100111111110100000010;
REG[4909] <= 32'b11111101000000001111101011110010;
REG[4910] <= 32'b11111001000000000000011100001001;
REG[4911] <= 32'b11101100111101011111110100011000;
REG[4912] <= 32'b00001011000001001111100011110100;
REG[4913] <= 32'b00000001111111101111111100000100;
REG[4914] <= 32'b11110000111111011111110011111010;
REG[4915] <= 32'b00000100000000011110101011111011;
REG[4916] <= 32'b00000010111111110000101100000110;
REG[4917] <= 32'b11110100111111001111100111111000;
REG[4918] <= 32'b11101010111110011111010111111101;
REG[4919] <= 32'b11110111111111001111010111110000;
REG[4920] <= 32'b11110110111110000000000011111001;
REG[4921] <= 32'b11110011111111000000010100000100;
REG[4922] <= 32'b00001001111110010000100000000000;
REG[4923] <= 32'b00000010111100010000001111110001;
REG[4924] <= 32'b00000011111110100000001000000100;
REG[4925] <= 32'b00000111111100101111111111111011;
REG[4926] <= 32'b00010010000010001111110111101100;
REG[4927] <= 32'b11110011111001011111010011110111;
REG[4928] <= 32'b00000100111100001111100011110011;
REG[4929] <= 32'b00000001111101001111011111111111;
REG[4930] <= 32'b00000100111001101111110111111011;
REG[4931] <= 32'b11111101000000001111010011110110;
REG[4932] <= 32'b11111011111110100000000000000110;
REG[4933] <= 32'b00000011111110111111011011111111;
REG[4934] <= 32'b00000111000010000000100011110101;
REG[4935] <= 32'b11110000111111011111101100001101;
REG[4936] <= 32'b11111110111100111111001100001001;
REG[4937] <= 32'b00000001000101110000100111110100;
REG[4938] <= 32'b11111011000101000000011000010111;
REG[4939] <= 32'b00000011111101111111111111111011;
REG[4940] <= 32'b00000101111101101110111111111111;
REG[4941] <= 32'b00000011111110100000000011110100;
REG[4942] <= 32'b11111001111111110000100111111000;
REG[4943] <= 32'b11111001111101001111110000000110;
REG[4944] <= 32'b00011010000001011111010111110101;
REG[4945] <= 32'b11110101111110010001111000011100;
REG[4946] <= 32'b00000100000001000000000011110000;
REG[4947] <= 32'b00011001000100011111100111110110;
REG[4948] <= 32'b00000000000000110000001000001111;
REG[4949] <= 32'b00011101000010010000100000001101;
REG[4950] <= 32'b11110101000001000001101100010000;
REG[4951] <= 32'b00010100000110111111111100001010;
REG[4952] <= 32'b00001110000001100000001000001000;
REG[4953] <= 32'b11111110111100100000000011110111;
REG[4954] <= 32'b11101010111110000001110000001011;
REG[4955] <= 32'b00000111111111011111011100000001;
REG[4956] <= 32'b11111000111100110000001011110001;
REG[4957] <= 32'b11110101111111011111010011101011;
REG[4958] <= 32'b11110000111111011110110000000110;
REG[4959] <= 32'b00000110000001000000100000000111;
REG[4960] <= 32'b11110110000010100000100111111111;
REG[4961] <= 32'b11110111111100111110010011101101;
REG[4962] <= 32'b11110011111101101111011000001010;
REG[4963] <= 32'b00000110111110111110111011101110;
REG[4964] <= 32'b11111110000001011111100011111110;
REG[4965] <= 32'b11101110111100101111011100000010;
REG[4966] <= 32'b11101001111011001111011100000000;
REG[4967] <= 32'b00000011000000001111111011111011;
REG[4968] <= 32'b00001000000100000001000011111110;
REG[4969] <= 32'b00000001111111010000100000010110;
REG[4970] <= 32'b00001001111111011111110011111000;
REG[4971] <= 32'b11110101111101010000001111111011;
REG[4972] <= 32'b11110000111101111111010111111000;
REG[4973] <= 32'b00000010000000011111101111111101;
REG[4974] <= 32'b11110000111101101111101011111100;
REG[4975] <= 32'b11110111111111111111001111111100;
REG[4976] <= 32'b00010111000100000000101100001000;
REG[4977] <= 32'b11110001111111010000001000000100;
REG[4978] <= 32'b00000110000001101110111011110011;
REG[4979] <= 32'b11110111111111111111110100000100;
REG[4980] <= 32'b00010101000011010000010000000001;
REG[4981] <= 32'b11110000000000100000010000001100;
REG[4982] <= 32'b00010010000101000000110100000011;
REG[4983] <= 32'b00000100000000110000000100000001;
REG[4984] <= 32'b11111101111110000000011100011100;
REG[4985] <= 32'b00000111000111111111111100010011;
REG[4986] <= 32'b11111000111101001111101000011000;
REG[4987] <= 32'b11110101000000010000011100000011;
REG[4988] <= 32'b00000010111111011111100111110000;
REG[4989] <= 32'b11111111000001101111001111110110;
REG[4990] <= 32'b11111111000001000000011100000010;
REG[4991] <= 32'b11110101111101100000000011101101;
REG[4992] <= 32'b00001001000001011111111111110011;
REG[4993] <= 32'b00010111111100011111111100000101;
REG[4994] <= 32'b00000100111101001111100011110101;
REG[4995] <= 32'b11110000000111000000101100000011;
REG[4996] <= 32'b11110001111110000000000000010001;
REG[4997] <= 32'b11110111000001011111111000000011;
REG[4998] <= 32'b11111010111111101111111000001011;
REG[4999] <= 32'b11111010111111111111101011111100;
REG[5000] <= 32'b00000000000010101111111111111010;
REG[5001] <= 32'b00000001111110011111110100000000;
REG[5002] <= 32'b11111000111110101111001100000010;
REG[5003] <= 32'b00001100111111010000111000000101;
REG[5004] <= 32'b00000001000010100000110000000110;
REG[5005] <= 32'b00001101000011110000010100001011;
REG[5006] <= 32'b00000111111111001111101000000110;
REG[5007] <= 32'b11111001111110011111110100000010;
REG[5008] <= 32'b11111111111101101111101100000100;
REG[5009] <= 32'b11111011111101111111000111110011;
REG[5010] <= 32'b00000001000001101111100111110010;
REG[5011] <= 32'b11110001111010101111001011111011;
REG[5012] <= 32'b00000011000001100000001011111101;
REG[5013] <= 32'b11110110111110111111010000001001;
REG[5014] <= 32'b11111101111101101111111100000110;
REG[5015] <= 32'b00000010000001000000010011111000;
REG[5016] <= 32'b00000110000000011110111000000010;
REG[5017] <= 32'b11101111111100100000110100010011;
REG[5018] <= 32'b11110110000001111110111100000010;
REG[5019] <= 32'b00000010000110010000011100000010;
REG[5020] <= 32'b11110000000101101110111111111111;
REG[5021] <= 32'b11111110111110101110111111101101;
REG[5022] <= 32'b00000100000011111111111111111110;
REG[5023] <= 32'b11111000111011110000100100000101;
REG[5024] <= 32'b00000001111101111111111011101100;
REG[5025] <= 32'b11101010000000111111111111110010;
REG[5026] <= 32'b11111000000010001111100000001110;
REG[5027] <= 32'b00001110111011111110111100000000;
REG[5028] <= 32'b11111101000010110001001111111101;
REG[5029] <= 32'b11110100111110001111001000000001;
REG[5030] <= 32'b00010010111110011111101111111100;
REG[5031] <= 32'b11111010111101010000001011111000;
REG[5032] <= 32'b11111010111111110000000111110101;
REG[5033] <= 32'b00000101111110001111100011111011;
REG[5034] <= 32'b00000000111111101111111011110101;
REG[5035] <= 32'b11111011111110010000011100000010;
REG[5036] <= 32'b11111100111101101111101000001110;
REG[5037] <= 32'b11111010111111001111110000000011;
REG[5038] <= 32'b11111001000100111111010111111010;
REG[5039] <= 32'b00010000111001011111011100100011;
REG[5040] <= 32'b00000111000110110001101011111001;
REG[5041] <= 32'b11111101000100001111101100000100;
REG[5042] <= 32'b00000101111110010000000011111011;
REG[5043] <= 32'b11111000000001101111011100001000;
REG[5044] <= 32'b00001111111110101111011100000101;
REG[5045] <= 32'b11111100111111010000100100000011;
REG[5046] <= 32'b11110101111111101111000000001111;
REG[5047] <= 32'b11111101111111000000111100001011;
REG[5048] <= 32'b00000010000000001111101011111001;
REG[5049] <= 32'b00001001000000111111100111111101;
REG[5050] <= 32'b00000000000000101111011111111100;
REG[5051] <= 32'b11111110000001000000011100001000;
REG[5052] <= 32'b11110101111111101111110000001100;
REG[5053] <= 32'b00110010001011111111000111111110;
REG[5054] <= 32'b00000100000111101111110011111100;
REG[5055] <= 32'b11111011000000111111110100000001;
REG[5056] <= 32'b11110001111110010000011100000011;
REG[5057] <= 32'b00000010000001001111101011110010;
REG[5058] <= 32'b11111111111110101111101011111111;
REG[5059] <= 32'b00001110111110111111011000000101;
REG[5060] <= 32'b00000011111111100000010111111000;
REG[5061] <= 32'b11110110111101001111010100001000;
REG[5062] <= 32'b11110110111111001111011011101011;
REG[5063] <= 32'b11111110000001001111001111110001;
REG[5064] <= 32'b11110100111100101111111011111101;
REG[5065] <= 32'b11111000111110100001101100000101;
REG[5066] <= 32'b00000010111011100000011000010010;
REG[5067] <= 32'b11110001111110110000001011101101;
REG[5068] <= 32'b00010001111100100001001000010000;
REG[5069] <= 32'b00000011111111000010111000001010;
REG[5070] <= 32'b00000001111111010000011011111001;
REG[5071] <= 32'b11110100000100010000111100011110;
REG[5072] <= 32'b00011011111101101110010100011001;
REG[5073] <= 32'b00000000000011110001010011110110;
REG[5074] <= 32'b00001011011001101111101011111010;
REG[5075] <= 32'b11101001111110001111101111111010;
REG[5076] <= 32'b11111100111110111110010111110101;
REG[5077] <= 32'b11111001111110110000000000010001;
REG[5078] <= 32'b11111101111010101111011111111100;
REG[5079] <= 32'b11111000111111110000001100000101;
REG[5080] <= 32'b00000000111100011111001011111111;
REG[5081] <= 32'b00001000000000111111100011110111;
REG[5082] <= 32'b00000100000001010000111000001001;
REG[5083] <= 32'b11110100111110100000100011111011;
REG[5084] <= 32'b11111100111101111111010111111010;
REG[5085] <= 32'b00010011000011011111111000000000;
REG[5086] <= 32'b00000000111101100000010111111110;
REG[5087] <= 32'b00000010111110011111100011110000;
REG[5088] <= 32'b11110110111101101111001000000001;
REG[5089] <= 32'b11111011111100101111110011111001;
REG[5090] <= 32'b11110100111110101111101111111011;
REG[5091] <= 32'b11110110111100101110110011111000;
REG[5092] <= 32'b11111100000000010000001100000000;
REG[5093] <= 32'b00000001111111010001100000000000;
REG[5094] <= 32'b00001000001000110001011111110011;
REG[5095] <= 32'b00000100111111110000000100000100;
REG[5096] <= 32'b00000001111101101111101111110010;
REG[5097] <= 32'b11110011111101001110011111110010;
REG[5098] <= 32'b00010000000000010000000100000011;
REG[5099] <= 32'b11110011111110000010011100001011;
REG[5100] <= 32'b00001000000010101111111000000010;
REG[5101] <= 32'b00000011111101010000001000000110;
REG[5102] <= 32'b11111111000100101111110011110010;
REG[5103] <= 32'b00011010000100110000011011101110;
REG[5104] <= 32'b11110101111101010001111000000001;
REG[5105] <= 32'b11111001000010010001011000011100;
REG[5106] <= 32'b11111011000010000000001011111000;
REG[5107] <= 32'b11110100111111001111100100001101;
REG[5108] <= 32'b00000000111101111110111111111111;
REG[5109] <= 32'b11111011000011010000001111110110;
REG[5110] <= 32'b11110111111111100000111000000011;
REG[5111] <= 32'b00000100111110101111111111111010;
REG[5112] <= 32'b00000001111110100000000111111011;
REG[5113] <= 32'b11111010111111010001010100001100;
REG[5114] <= 32'b00000001111110111111010011110011;
REG[5115] <= 32'b00000010000000011111110000000101;
REG[5116] <= 32'b00000000111110010000000011111101;
REG[5117] <= 32'b11111110111111111111111111111101;
REG[5118] <= 32'b11111110000000011111101111110100;
REG[5119] <= 32'b11110000111100100000001000000010;
REG[5120] <= 32'b00000011111101111111011111110110;
REG[5121] <= 32'b11110111111101001111000111110001;
REG[5122] <= 32'b11111100111110100000111100001000;
REG[5123] <= 32'b11111110111011101111010111111010;
REG[5124] <= 32'b00000111000001110000010000101000;
REG[5125] <= 32'b00011001111111001111110011111011;
REG[5126] <= 32'b00000011000110110000011100000101;
REG[5127] <= 32'b11111010111111111111111111110111;
REG[5128] <= 32'b11101011111111101111111011111110;
REG[5129] <= 32'b11111101111101100000011100001000;
REG[5130] <= 32'b00000111000101010000001100000010;
REG[5131] <= 32'b11111000000000001111110100000101;
REG[5132] <= 32'b00000100111111011111111111111101;
REG[5133] <= 32'b11111110000001100000010100010010;
REG[5134] <= 32'b11111000111101110000001111111011;
REG[5135] <= 32'b00000110000010011111000111111110;
REG[5136] <= 32'b00001010111111011111110011111011;
REG[5137] <= 32'b11111001000100010000010100000100;
REG[5138] <= 32'b11111111111101100000111000010101;
REG[5139] <= 32'b00000001111111001111110011110110;
REG[5140] <= 32'b00010010000100110001001000001010;
REG[5141] <= 32'b00001001000000011111111100000011;
REG[5142] <= 32'b11110110111100101110111100010110;
REG[5143] <= 32'b00001111000010001110111111110110;
REG[5144] <= 32'b11111011000011010000101000000001;
REG[5145] <= 32'b00000010111110001111101111110111;
REG[5146] <= 32'b00000010000000000000000100000001;
REG[5147] <= 32'b00000001000010000000010111111110;
REG[5148] <= 32'b00000010000010110000100100000100;
REG[5149] <= 32'b11111100111111001111110000000001;
REG[5150] <= 32'b11111010000010010000001011111001;
REG[5151] <= 32'b11110111111110010000001111110111;
REG[5152] <= 32'b11111010111111001111101111111001;
REG[5153] <= 32'b00000001111100111111101111111100;
REG[5154] <= 32'b00000001000001110000110011110001;
REG[5155] <= 32'b11111110000010000000100100001010;
REG[5156] <= 32'b00000110111111011111101011110111;
REG[5157] <= 32'b00001011000010010000001111111100;
REG[5158] <= 32'b11110100111110000000010100000101;
REG[5159] <= 32'b00000000000000000000000011111011;
REG[5160] <= 32'b11111001111101001110111100010111;
REG[5161] <= 32'b11110001111011100000110100101010;
REG[5162] <= 32'b11111001000110101111001011110001;
REG[5163] <= 32'b00010101001101110000100100010001;
REG[5164] <= 32'b00000010111110000000000100000011;
REG[5165] <= 32'b00000001111110011111010111110001;
REG[5166] <= 32'b00001001000011000001001011110000;
REG[5167] <= 32'b11101101111100100000101000010001;
REG[5168] <= 32'b00001010000100110000110100000010;
REG[5169] <= 32'b11111000000000101111111011110001;
REG[5170] <= 32'b11101100000000101111111111111111;
REG[5171] <= 32'b00000001111011001110100100000110;
REG[5172] <= 32'b11110101111100011111100011111001;
REG[5173] <= 32'b11111010000010101111111000000001;
REG[5174] <= 32'b00000000000000010000001111110011;
REG[5175] <= 32'b00001111000011100000110111111101;
REG[5176] <= 32'b11111011111111001111111000000000;
REG[5177] <= 32'b00000000000010110000011100010010;
REG[5178] <= 32'b00001100000000001111101000010010;
REG[5179] <= 32'b00000010000110100000010011110101;
REG[5180] <= 32'b11101110000000001111110100001100;
REG[5181] <= 32'b11110101111110111111111011111001;
REG[5182] <= 32'b00000011111111000000010000000100;
REG[5183] <= 32'b00000001111110100000111000000001;
REG[5184] <= 32'b00010101000110110001010111110111;
REG[5185] <= 32'b11111101111111000000010100001110;
REG[5186] <= 32'b00000100000010100000011011111010;
REG[5187] <= 32'b00000011000000010000010100001101;
REG[5188] <= 32'b11110101000000100000000011111001;
REG[5189] <= 32'b11111110000010011111010100000001;
REG[5190] <= 32'b11111111111100101111100000001011;
REG[5191] <= 32'b11110111000000111111111000000111;
REG[5192] <= 32'b00000101111111000010000000011101;
REG[5193] <= 32'b11110111111110011111010100000100;
REG[5194] <= 32'b00001100111111110000010100001100;
REG[5195] <= 32'b00010011111110011111110111111000;
REG[5196] <= 32'b11111011000000000000000011111010;
REG[5197] <= 32'b11111111000001101111111000100100;
REG[5198] <= 32'b11111011111101001111011000000011;
REG[5199] <= 32'b11110111000111000000101011100111;
REG[5200] <= 32'b00000101111111000000000100001001;
REG[5201] <= 32'b00000010000010110001011100000111;
REG[5202] <= 32'b11101110111010011110110011111101;
REG[5203] <= 32'b00000110000001110000001100000011;
REG[5204] <= 32'b00001000111110111111101111111110;
REG[5205] <= 32'b11111100111111001111001111110101;
REG[5206] <= 32'b00100101111111000000100000001110;
REG[5207] <= 32'b11111100111110110001110111110000;
REG[5208] <= 32'b00010110001000001111110011110101;
REG[5209] <= 32'b00010000000001000000011100000110;
REG[5210] <= 32'b00000010000100010000010111110111;
REG[5211] <= 32'b00010100000011110000011100001000;
REG[5212] <= 32'b00000111111101000000110100000111;
REG[5213] <= 32'b11111110111101111111110011111000;
REG[5214] <= 32'b11111101111110101111100111101110;
REG[5215] <= 32'b11100110111100001111011111111000;
REG[5216] <= 32'b11111001111010111110001011101101;
REG[5217] <= 32'b11111100111110010000100100000010;
REG[5218] <= 32'b11110101111111001111110111111111;
REG[5219] <= 32'b00000000111110001111011000001000;
REG[5220] <= 32'b00001100000010110000100111110101;
REG[5221] <= 32'b11101111111001110000001000000110;
REG[5222] <= 32'b00001100000001110000100011101110;
REG[5223] <= 32'b11111000111110101110111011111111;
REG[5224] <= 32'b11110110111101010000001000000101;
REG[5225] <= 32'b11111100000001001111101000000010;
REG[5226] <= 32'b00000010111111001111110000000101;
REG[5227] <= 32'b11110101111111010000100100001010;
REG[5228] <= 32'b00000110111110110000001100001000;
REG[5229] <= 32'b11111011111111111111101100000001;
REG[5230] <= 32'b11110110111101100000010000000001;
REG[5231] <= 32'b11111010111101111111000111110001;
REG[5232] <= 32'b11111001000001111111101000000011;
REG[5233] <= 32'b00000010111100101111011000001110;
REG[5234] <= 32'b11111001000010110000000111111011;
REG[5235] <= 32'b11110111111110101110100000001111;
REG[5236] <= 32'b11111111111101111111110100001000;
REG[5237] <= 32'b00001100111111100000011011101110;
REG[5238] <= 32'b00000011000001101111101000000001;
REG[5239] <= 32'b00000100111010110000001111111001;
REG[5240] <= 32'b11111110000001000000001111101110;
REG[5241] <= 32'b11110001111110000000101100001101;
REG[5242] <= 32'b00001011000100001111010111110110;
REG[5243] <= 32'b00001011000000000000010000001110;
REG[5244] <= 32'b11101001111101000000010011110111;
REG[5245] <= 32'b11110100000001111110111000000011;
REG[5246] <= 32'b00001101111110100000001011111000;
REG[5247] <= 32'b11100000000001000001010011111010;
REG[5248] <= 32'b11111101000001011110111011110101;
REG[5249] <= 32'b00001101000000100001001000000110;
REG[5250] <= 32'b11111100111110111111100000000010;
REG[5251] <= 32'b11110010111111110000001011111110;
REG[5252] <= 32'b11111101000010001111000011101011;
REG[5253] <= 32'b11111100111110001111110000000100;
REG[5254] <= 32'b11110010111100000000011000000001;
REG[5255] <= 32'b11111111111011111111101111110100;
REG[5256] <= 32'b00100101000011011111100000000010;
REG[5257] <= 32'b00001011000001100001111000001110;
REG[5258] <= 32'b00000001000001100000000000000101;
REG[5259] <= 32'b00000111000000000000000000000101;
REG[5260] <= 32'b11111101000011001111111111110110;
REG[5261] <= 32'b11110011111110001111011111111010;
REG[5262] <= 32'b00000010000010110000010000000100;
REG[5263] <= 32'b11110110111011110000110100010001;
REG[5264] <= 32'b00000001111111010000100100010101;
REG[5265] <= 32'b00010011000010010000000000000010;
REG[5266] <= 32'b00000101000001110000110011111101;
REG[5267] <= 32'b11111011000000011111101000001000;
REG[5268] <= 32'b00001111000011011111100000000101;
REG[5269] <= 32'b00001101111111000001000111111000;
REG[5270] <= 32'b11101010111110111111100111110011;
REG[5271] <= 32'b00000010111110111101111100000110;
REG[5272] <= 32'b11111011000000101111110011110010;
REG[5273] <= 32'b00000101111111111111100011110100;
REG[5274] <= 32'b11110111111110000000001111111100;
REG[5275] <= 32'b11110000111100111111101111110000;
REG[5276] <= 32'b00000010111101111111010011111110;
REG[5277] <= 32'b11111110111111011111000011110010;
REG[5278] <= 32'b00001010000111011111101011111111;
REG[5279] <= 32'b11110101111101110000100000011011;
REG[5280] <= 32'b11110100111111001111010100000011;
REG[5281] <= 32'b11111010000001110000011000001001;
REG[5282] <= 32'b00000110111110101111110100001000;
REG[5283] <= 32'b11111111000000110000100011110001;
REG[5284] <= 32'b11110110111110000000111000000100;
REG[5285] <= 32'b11111100111100101111010011111011;
REG[5286] <= 32'b11101111000011000000111011101001;
REG[5287] <= 32'b11111001000000111101101100011110;
REG[5288] <= 32'b00100011111010101111101000000100;
REG[5289] <= 32'b11101110000011100001011011101100;
REG[5290] <= 32'b11111001000001010000100011110011;
REG[5291] <= 32'b11110100000100110010010000000001;
REG[5292] <= 32'b00011011111110011111011100001010;
REG[5293] <= 32'b00100100000011100001000000001000;
REG[5294] <= 32'b00000010000010110000110100010000;
REG[5295] <= 32'b11101110111011101111001011111101;
REG[5296] <= 32'b11111111111111001110111011110010;
REG[5297] <= 32'b11110011111111001111010011111110;
REG[5298] <= 32'b11110011111101011111101100001010;
REG[5299] <= 32'b00000100000000010000001000000010;
REG[5300] <= 32'b00001100111110101111111011101110;
REG[5301] <= 32'b00010101111101111111000111111000;
REG[5302] <= 32'b11111110111111010000000011101100;
REG[5303] <= 32'b00000001111101110000001111111001;
REG[5304] <= 32'b00000010000010110001010011111111;
REG[5305] <= 32'b11111010000001101111111011111100;
REG[5306] <= 32'b00010000000000001110111000011100;
REG[5307] <= 32'b11111010111100110000000000000110;
REG[5308] <= 32'b11110001111111100000001111111111;
REG[5309] <= 32'b00000001111101111111010111110011;
REG[5310] <= 32'b00001111111111110000011100000101;
REG[5311] <= 32'b00000101111101010000110111111111;
REG[5312] <= 32'b00000100000011010000010000001000;
REG[5313] <= 32'b11110111111101011111001011111010;
REG[5314] <= 32'b11111011000000001110111111101111;
REG[5315] <= 32'b11101011111110111110110011101101;
REG[5316] <= 32'b00000000000010101111111111111011;
REG[5317] <= 32'b00000000000000000000000000000011;
REG[5318] <= 32'b00000011111011111111000111111100;
REG[5319] <= 32'b00001001111101101111111011111100;
REG[5320] <= 32'b11111101111110010000111111110110;
REG[5321] <= 32'b00000101111101001111110111110110;
REG[5322] <= 32'b11110111000010010000011100000001;
REG[5323] <= 32'b11111000111110001111011011111001;
REG[5324] <= 32'b11110110111111111111010111110101;
REG[5325] <= 32'b00001000111111111110101111111010;
REG[5326] <= 32'b11110001000000000000010100000000;
REG[5327] <= 32'b00000111000000011111011111111011;
REG[5328] <= 32'b00011001000010000000011100000010;
REG[5329] <= 32'b00000001111110110000000000000010;
REG[5330] <= 32'b00000111000000111111111111111110;
REG[5331] <= 32'b00000100000000010001010011111101;
REG[5332] <= 32'b00001100000000000000000000000010;
REG[5333] <= 32'b00010011000001001111111000000000;
REG[5334] <= 32'b11110011111110010000011100000111;
REG[5335] <= 32'b00010001000011001110101111111100;
REG[5336] <= 32'b00000001111100001111011111111111;
REG[5337] <= 32'b11110110111111001111110111110011;
REG[5338] <= 32'b11111011111101111111001011111011;
REG[5339] <= 32'b11111010111010001111011011110110;
REG[5340] <= 32'b11111010111110011111101111101111;
REG[5341] <= 32'b11100000111101101111101111110100;
REG[5342] <= 32'b11110011111100111111001100001010;
REG[5343] <= 32'b11110010111101001111011011111101;
REG[5344] <= 32'b00000000111101101111101000000110;
REG[5345] <= 32'b00001010000000110000000011111010;
REG[5346] <= 32'b00000110000001110000011100001101;
REG[5347] <= 32'b00010010111111000000000100001101;
REG[5348] <= 32'b00010000000011001111110111111001;
REG[5349] <= 32'b11110101111100000000111011100111;
REG[5350] <= 32'b11110001111110011111101111101111;
REG[5351] <= 32'b11111011111011111111110111111100;
REG[5352] <= 32'b00000000111101011111101111110101;
REG[5353] <= 32'b00001010000010100000000000000000;
REG[5354] <= 32'b00000110111111000000001000001001;
REG[5355] <= 32'b11110101111111110000110100000000;
REG[5356] <= 32'b00000011000000001111001111111101;
REG[5357] <= 32'b00001111000000011111111111111010;
REG[5358] <= 32'b11101010111010111111010100000001;
REG[5359] <= 32'b11110110000010101111000111101001;
REG[5360] <= 32'b11101101111101101101110111110111;
REG[5361] <= 32'b11110100111011111111011111111010;
REG[5362] <= 32'b11110000000001000000100111111001;
REG[5363] <= 32'b11111000000010010000110000001000;
REG[5364] <= 32'b00000100000001000000100100001011;
REG[5365] <= 32'b00000011000100001111100011111110;
REG[5366] <= 32'b11111010000011110000100000001101;
REG[5367] <= 32'b11110101111100111111110100001100;
REG[5368] <= 32'b11110010111100101111100111101111;
REG[5369] <= 32'b11111010000100011111010011110000;
REG[5370] <= 32'b11111011111101100000001000010000;
REG[5371] <= 32'b11111100111110001111001111111101;
REG[5372] <= 32'b00000001111111110000011100000001;
REG[5373] <= 32'b11111001111111100000010111111001;
REG[5374] <= 32'b00010001000000101111101000000000;
REG[5375] <= 32'b00001101111111110000100000000001;
REG[5376] <= 32'b11101111111110001111110011111010;
REG[5377] <= 32'b11110100111110101110101011101101;
REG[5378] <= 32'b11101100111111010000000000000011;
REG[5379] <= 32'b11101010111011001110111011111111;
REG[5380] <= 32'b00001000000010011110110111101001;
REG[5381] <= 32'b11110101111101011110110111101110;
REG[5382] <= 32'b11111101111001101110110011111001;
REG[5383] <= 32'b11110111111100100000011111101100;
REG[5384] <= 32'b11101110111110011111011111110110;
REG[5385] <= 32'b11110010111100111111100011111101;
REG[5386] <= 32'b00000000000001011111100011111001;
REG[5387] <= 32'b00000111111101100000100100000000;
REG[5388] <= 32'b11110100111010001111111100010010;
REG[5389] <= 32'b00101010111110001111101000000011;
REG[5390] <= 32'b00000100111111111111111100001001;
REG[5391] <= 32'b00001011111111011111000000000110;
REG[5392] <= 32'b11111000111100110001011100000000;
REG[5393] <= 32'b11111111111110100000010100001101;
REG[5394] <= 32'b11110101111100001110111000000111;
REG[5395] <= 32'b00011010000000010000100000000001;
REG[5396] <= 32'b11110010111110000000100111110010;
REG[5397] <= 32'b00010100000010011111001011111101;
REG[5398] <= 32'b11111110000000011111101011111011;
REG[5399] <= 32'b11111111000001111111001011110000;
REG[5400] <= 32'b11110101111100001111111000010110;
REG[5401] <= 32'b00000100111110101111101111111011;
REG[5402] <= 32'b11111101000101110001000000001011;
REG[5403] <= 32'b11110110111110011111101100001001;
REG[5404] <= 32'b11111110111101001111010111111000;
REG[5405] <= 32'b11111100000011000000110011111011;
REG[5406] <= 32'b11110011111011101111000100000000;
REG[5407] <= 32'b11111101111100001111100100000000;
REG[5408] <= 32'b11111111000010101111001111110110;
REG[5409] <= 32'b11101111000000010000101100000011;
REG[5410] <= 32'b11110100111101111110111111110010;
REG[5411] <= 32'b00000100111111111111011111111001;
REG[5412] <= 32'b11110110111011111111001011110110;
REG[5413] <= 32'b11111000111100110000101011111100;
REG[5414] <= 32'b11110110000000100001110000010010;
REG[5415] <= 32'b11110010111010101110111000000101;
REG[5416] <= 32'b00011001000100010000100000010000;
REG[5417] <= 32'b00001000001000101111111111110110;
REG[5418] <= 32'b11101111000001100000100000001010;
REG[5419] <= 32'b11110010111101010000011100001001;
REG[5420] <= 32'b11111100111001011111010111110100;
REG[5421] <= 32'b00000011111100011111101111111101;
REG[5422] <= 32'b11111010111100100001001011110111;
REG[5423] <= 32'b11111000111111100000001011111100;
REG[5424] <= 32'b00000110000000001111000100001101;
REG[5425] <= 32'b00011001001010111111111000010110;
REG[5426] <= 32'b00001011000100111111100111111101;
REG[5427] <= 32'b00000011111110010001010000011010;
REG[5428] <= 32'b11110000111110011111000111100110;
REG[5429] <= 32'b00001101000001011111101000000100;
REG[5430] <= 32'b00001101000000101111111000010101;
REG[5431] <= 32'b00010001000011000000110000000101;
REG[5432] <= 32'b11111111000001000000000011111000;
REG[5433] <= 32'b00000101000000100000010000000011;
REG[5434] <= 32'b00001011000000010000000011110100;
REG[5435] <= 32'b11111110111100101111001000001001;
REG[5436] <= 32'b00011101111011011111001011110110;
REG[5437] <= 32'b11110100000100100001001111110010;
REG[5438] <= 32'b11110010111010001111010000001110;
REG[5439] <= 32'b00000110000000010000001100010000;
REG[5440] <= 32'b00000001111110100000110100000000;
REG[5441] <= 32'b11111100000100100000010011110001;
REG[5442] <= 32'b00001011000000111111111000010000;
REG[5443] <= 32'b00000110111111001111100100001000;
REG[5444] <= 32'b00010001111101011111010000000101;
REG[5445] <= 32'b00000100111101100000010011101100;
REG[5446] <= 32'b11110000000001100000000100001000;
REG[5447] <= 32'b00000111111110100000110000001110;
REG[5448] <= 32'b00000101111101001110111011110011;
REG[5449] <= 32'b00000111000000000000110011110110;
REG[5450] <= 32'b11111111111100110000011011111111;
REG[5451] <= 32'b00001101111011010000001000001011;
REG[5452] <= 32'b00001001000011111111011111111110;
REG[5453] <= 32'b00001011000100001110110111110000;
REG[5454] <= 32'b11111010111101101111101100001110;
REG[5455] <= 32'b11110010000000000000101011110000;
REG[5456] <= 32'b11110001111111101111110000001001;
REG[5457] <= 32'b11101110111110011111100111111000;
REG[5458] <= 32'b11110001111111101111100111111011;
REG[5459] <= 32'b11111000111101101111001100000000;
REG[5460] <= 32'b00000100111110111111010100000111;
REG[5461] <= 32'b00001001000000110000000111111001;
REG[5462] <= 32'b11111100111111011111100011111111;
REG[5463] <= 32'b00010101000001110000010111110101;
REG[5464] <= 32'b11111011111110100001111000001000;
REG[5465] <= 32'b00001010111110011111111011110110;
REG[5466] <= 32'b11111001111111110000100011111001;
REG[5467] <= 32'b00010011000000110000000111110111;
REG[5468] <= 32'b00000000111101010000011111111100;
REG[5469] <= 32'b00000101111110001111011011111110;
REG[5470] <= 32'b11111101111101011111011011111011;
REG[5471] <= 32'b11111110000100010000001100000100;
REG[5472] <= 32'b11101110111010001111000100000000;
REG[5473] <= 32'b00000010000000111111100011110101;
REG[5474] <= 32'b11110010111111011111011011111011;
REG[5475] <= 32'b11110000111101100001010000001000;
REG[5476] <= 32'b00000001111110011111011111110010;
REG[5477] <= 32'b00001011111111101111111011111010;
REG[5478] <= 32'b11111000111011010000101011111010;
REG[5479] <= 32'b11111000111111111111110000000010;
REG[5480] <= 32'b00000110111010101110100100001111;
REG[5481] <= 32'b11110111000001000000010111111001;
REG[5482] <= 32'b11101011000100001111100111111010;
REG[5483] <= 32'b00000000000000110000010000100101;
REG[5484] <= 32'b11111111000010110000100011111111;
REG[5485] <= 32'b00000011111110010000011100000000;
REG[5486] <= 32'b11111011111101101110111111111101;
REG[5487] <= 32'b00001100111111001111010111110110;
REG[5488] <= 32'b11110100111111000000010000001000;
REG[5489] <= 32'b00010011000001110000011100000000;
REG[5490] <= 32'b11111101000001110001000011110010;
REG[5491] <= 32'b11110000111111011111010111111011;
REG[5492] <= 32'b11111111111110010000000000000100;
REG[5493] <= 32'b00000101000000100000010000001100;
REG[5494] <= 32'b00000100111110011111101011110111;
REG[5495] <= 32'b00000000000000000000110100000010;
REG[5496] <= 32'b00001101111110110000000111110110;
REG[5497] <= 32'b11111000111101000000001111111101;
REG[5498] <= 32'b00001010111101001110111000001010;
REG[5499] <= 32'b11110101111011000000000111111010;
REG[5500] <= 32'b11111110000010011111111000000000;
REG[5501] <= 32'b00000010000010110000000100001100;
REG[5502] <= 32'b00001001000011011111100100001001;
REG[5503] <= 32'b00000100000001110000011011111001;
REG[5504] <= 32'b11111101000001000000100011110110;
REG[5505] <= 32'b00000000111111011111101000001101;
REG[5506] <= 32'b00010011111111101111111111110111;
REG[5507] <= 32'b11111100111110101111111011111010;
REG[5508] <= 32'b11111010111110011111111011110000;
REG[5509] <= 32'b11111001111110011111111111110110;
REG[5510] <= 32'b11110110000000011111110011111100;
REG[5511] <= 32'b11111101111101111111001000000000;
REG[5512] <= 32'b11111001111110100000101111111011;
REG[5513] <= 32'b11110011111110101111011011111000;
REG[5514] <= 32'b00010100000010101111010111111110;
REG[5515] <= 32'b11110110111111000000000111111001;
REG[5516] <= 32'b11111001111100011111001000001010;
REG[5517] <= 32'b11110100111111000000011011110101;
REG[5518] <= 32'b11111101000100100000000000000111;
REG[5519] <= 32'b11111111000000110000110100001111;
REG[5520] <= 32'b00000000111111011111000011111111;
REG[5521] <= 32'b11111001000000101111100111111111;
REG[5522] <= 32'b11110011000000001110100111111101;
REG[5523] <= 32'b00000010000000000000010000000011;
REG[5524] <= 32'b11110001111110110000100000000011;
REG[5525] <= 32'b11110110111110011111011111111011;
REG[5526] <= 32'b00000011000001000000001011111010;
REG[5527] <= 32'b11111101111111011111111100000001;
REG[5528] <= 32'b00000001111110011111111000000000;
REG[5529] <= 32'b11110100000001011111100000000110;
REG[5530] <= 32'b00001010000011011111111000010110;
REG[5531] <= 32'b00001010000001101111110000000100;
REG[5532] <= 32'b11110101111101111111110011111111;
REG[5533] <= 32'b11111111000100100000100011111101;
REG[5534] <= 32'b11110101111011011111101100001110;
REG[5535] <= 32'b00000100111110111110111111110010;
REG[5536] <= 32'b11110110111101110000110100000001;
REG[5537] <= 32'b11111101000001000000011100001000;
REG[5538] <= 32'b00000010111110011110011011111001;
REG[5539] <= 32'b00000001000001011111110111110101;
REG[5540] <= 32'b11110000000001111111111100000010;
REG[5541] <= 32'b11110010111100101111000000010010;
REG[5542] <= 32'b00000111000000101111010111110011;
REG[5543] <= 32'b11110111000110001111111011111101;
REG[5544] <= 32'b11110010111100111111110011111110;
REG[5545] <= 32'b11110000111110101111011011110011;
REG[5546] <= 32'b11110111111101101111010111110001;
REG[5547] <= 32'b11111111000001110001000100000011;
REG[5548] <= 32'b00001001000010100000101011111101;
REG[5549] <= 32'b00000101000010101111111000001111;
REG[5550] <= 32'b00000011111110011111100100000010;
REG[5551] <= 32'b00000001000010100000010000001101;
REG[5552] <= 32'b00001001111100011111101100000100;
REG[5553] <= 32'b00001110000110000000111011111101;
REG[5554] <= 32'b00000000000010101111111100000100;
REG[5555] <= 32'b00000001000001000000010000001100;
REG[5556] <= 32'b11111000111100011111000000001001;
REG[5557] <= 32'b11110110000010101110101111110100;
REG[5558] <= 32'b11111101111100101111000011111000;
REG[5559] <= 32'b00000001000000010001010100000110;
REG[5560] <= 32'b11110001111101001111101111111001;
REG[5561] <= 32'b00001101000000000000001100011101;
REG[5562] <= 32'b11111101111111000000111111101110;
REG[5563] <= 32'b11100110111011101111111100000111;
REG[5564] <= 32'b00001100111110001111101100000000;
REG[5565] <= 32'b11111110111111001111110111111110;
REG[5566] <= 32'b11111101111110100000001111111001;
REG[5567] <= 32'b00000100000000011111100011110101;
REG[5568] <= 32'b11110111111101100000000100000111;
REG[5569] <= 32'b00000111111101010000000111111001;
REG[5570] <= 32'b11110010000001101111110000000001;
REG[5571] <= 32'b00000011000000110000000011100100;
REG[5572] <= 32'b11101101111110000000001100001100;
REG[5573] <= 32'b00001011111101100000001100000100;
REG[5574] <= 32'b11111100000100110001111111111100;
REG[5575] <= 32'b11101011000000111111110100000100;
REG[5576] <= 32'b00011101000010011111000100000110;
REG[5577] <= 32'b00001000000001100001101100010110;
REG[5578] <= 32'b11111011000010110000010000000000;
REG[5579] <= 32'b00000000111110111111001011111010;
REG[5580] <= 32'b11111101111110101111011011111100;
REG[5581] <= 32'b00001001000001011111011011101101;
REG[5582] <= 32'b11110001111110010000100000000101;
REG[5583] <= 32'b11111100111110011110100000001110;
REG[5584] <= 32'b00000101111111111111101011111000;
REG[5585] <= 32'b11101111000011011111011011111010;
REG[5586] <= 32'b11110010111101101110110100011110;
REG[5587] <= 32'b00010111000101000000000111110011;
REG[5588] <= 32'b11110110111011011110010111110001;
REG[5589] <= 32'b00001001111111111111100011110011;
REG[5590] <= 32'b11110110000010000000010111111111;
REG[5591] <= 32'b11111100000010001111011100000100;
REG[5592] <= 32'b11111100111110011111010100000010;
REG[5593] <= 32'b11110110111101011111111100000101;
REG[5594] <= 32'b00000010111110001111001111111000;
REG[5595] <= 32'b11111000111111001111001011111100;
REG[5596] <= 32'b11111110111101100000011011111010;
REG[5597] <= 32'b11111100000011110000010111110111;
REG[5598] <= 32'b00001010111110101111010111110100;
REG[5599] <= 32'b11110111111110011111110011111010;
REG[5600] <= 32'b11110100000000101111111000000110;
REG[5601] <= 32'b00000010111110000000001011111000;
REG[5602] <= 32'b00000001000101001111100011101110;
REG[5603] <= 32'b11111011111111001111101100000100;
REG[5604] <= 32'b11111100111101100000000100001010;
REG[5605] <= 32'b00000000111111100000111100000110;
REG[5606] <= 32'b00000100000011100000000100000100;
REG[5607] <= 32'b11111110111110111111101011110010;
REG[5608] <= 32'b11111000000000001111100011111010;
REG[5609] <= 32'b11111010111101010000000111111101;
REG[5610] <= 32'b00000100111111101111111111110111;
REG[5611] <= 32'b11111001111111111111111111111110;
REG[5612] <= 32'b11111110111010101111000011101111;
REG[5613] <= 32'b00000001000000011111111011111000;
REG[5614] <= 32'b11111011111100110000000000001011;
REG[5615] <= 32'b11110011000101110000001011101101;
REG[5616] <= 32'b00001000000010101111001111111001;
REG[5617] <= 32'b11111000111110010000001000000100;
REG[5618] <= 32'b11110111111111101111110111111000;
REG[5619] <= 32'b00011001000100100000000111110111;
REG[5620] <= 32'b11110111000000010000001111111011;
REG[5621] <= 32'b11111001000000111111011011111000;
REG[5622] <= 32'b00001010000000101111100011111101;
REG[5623] <= 32'b11111000000001001111100111110110;
REG[5624] <= 32'b11110110111010101111000111111001;
REG[5625] <= 32'b11111100000001000000010011101010;
REG[5626] <= 32'b11110010111111011111001011110100;
REG[5627] <= 32'b11111100111110001111111000010110;
REG[5628] <= 32'b00000001111100010000000100000011;
REG[5629] <= 32'b11101101000010101111100111110100;
REG[5630] <= 32'b00000110000000111111000100000111;
REG[5631] <= 32'b11111101111101111111001111111011;
REG[5632] <= 32'b11110011000010101111111100001010;
REG[5633] <= 32'b00000000111010101110110000001001;
REG[5634] <= 32'b00000001000010110000100011101011;
REG[5635] <= 32'b11111110000001111111010000001100;
REG[5636] <= 32'b00000010000010100001100100010000;
REG[5637] <= 32'b11111001000010101111110000000101;
REG[5638] <= 32'b00000011000010100000011000011010;
REG[5639] <= 32'b11111000111101110000000100000101;
REG[5640] <= 32'b00000001001011011111101011111000;
REG[5641] <= 32'b11110111000000111110110011110100;
REG[5642] <= 32'b11111011111010101110011111110111;
REG[5643] <= 32'b00000110111110111111100111110010;
REG[5644] <= 32'b11110100111111110001011000001001;
REG[5645] <= 32'b11110111000001001111110111111110;
REG[5646] <= 32'b11111101000000100000100111111110;
REG[5647] <= 32'b00001011000001011111101111111111;
REG[5648] <= 32'b11111000111100101111011111111101;
REG[5649] <= 32'b00001000000010100001010011101111;
REG[5650] <= 32'b11111110000010101111111111111111;
REG[5651] <= 32'b00000000111111011111111111101011;
REG[5652] <= 32'b11111100111110001111110100000111;
REG[5653] <= 32'b11111111111100111111101111111001;
REG[5654] <= 32'b00000000000001010000000100000001;
REG[5655] <= 32'b00001010000010110001001111111000;
REG[5656] <= 32'b00000111111100110000100000001000;
REG[5657] <= 32'b00001110111100000000000111110111;
REG[5658] <= 32'b00000001000010100000110111101111;
REG[5659] <= 32'b00000011111110011111110011110100;
REG[5660] <= 32'b11110110111111001110100011101101;
REG[5661] <= 32'b11111011111101001111100111110111;
REG[5662] <= 32'b11110010111100100000010011101110;
REG[5663] <= 32'b11110011111111011111011011110011;
REG[5664] <= 32'b11111010111101101111001011110011;
REG[5665] <= 32'b11111110111111011111101111110100;
REG[5666] <= 32'b11101100111100100000011011111101;
REG[5667] <= 32'b11110100111100101111001011110101;
REG[5668] <= 32'b11111110111110111110110111110111;
REG[5669] <= 32'b11111001000011001111111111110011;
REG[5670] <= 32'b11110011111101111111011111111110;
REG[5671] <= 32'b00001111000001011111111111111100;
REG[5672] <= 32'b11111101111011010000010011110111;
REG[5673] <= 32'b11101111000010010000000000000011;
REG[5674] <= 32'b11111101000110000001100100100101;
REG[5675] <= 32'b11110010000011010000011000011011;
REG[5676] <= 32'b00000010000011111110110100000110;
REG[5677] <= 32'b11111011000100011111011000000100;
REG[5678] <= 32'b00000100001000000000010100000011;
REG[5679] <= 32'b11111001000000001111011111110111;
REG[5680] <= 32'b11101101111100011111011000000100;
REG[5681] <= 32'b11110111111011100000000100001001;
REG[5682] <= 32'b00000110000000101111011000000000;
REG[5683] <= 32'b00000100000101100000001011110110;
REG[5684] <= 32'b11111100111111100000011000010011;
REG[5685] <= 32'b00001010111111000000010011111100;
REG[5686] <= 32'b11111110000101101111111000000110;
REG[5687] <= 32'b00010010111110101111111011110110;
REG[5688] <= 32'b11111100000011010001001011110011;
REG[5689] <= 32'b11111101111111111111011000000011;
REG[5690] <= 32'b11111100111111100000110000010110;
REG[5691] <= 32'b11111000000001100000111111111011;
REG[5692] <= 32'b11111110000010101111101011111111;
REG[5693] <= 32'b00001100111101111111011000000000;
REG[5694] <= 32'b00000000000010010000010000000001;
REG[5695] <= 32'b11111011000000001111111011111001;
REG[5696] <= 32'b11111011111100001110100011111001;
REG[5697] <= 32'b00000111111110001111100111110101;
REG[5698] <= 32'b11110001111101101111110111111101;
REG[5699] <= 32'b11111100000000011111001111110110;
REG[5700] <= 32'b11111110111110100001001011101100;
REG[5701] <= 32'b11110001000001101111100111111100;
REG[5702] <= 32'b00001110111011001111001000000101;
REG[5703] <= 32'b11110111111110100000100100000110;
REG[5704] <= 32'b00000001000100000000000111111010;
REG[5705] <= 32'b11110100000010110010001111111000;
REG[5706] <= 32'b00000100111101111111011011111001;
REG[5707] <= 32'b11111010111111110000000100000101;
REG[5708] <= 32'b00000011111011011110100000001101;
REG[5709] <= 32'b11111010111101101111011011111011;
REG[5710] <= 32'b11111010000010100000001100001101;
REG[5711] <= 32'b00000011111101001111010000000111;
REG[5712] <= 32'b00001111000011100000011011111010;
REG[5713] <= 32'b11111001000100001111111011111000;
REG[5714] <= 32'b11101101000000011111010111101011;
REG[5715] <= 32'b00000000000001111111001011111111;
REG[5716] <= 32'b11111111111101001111111000000000;
REG[5717] <= 32'b11111010000001111111100011111011;
REG[5718] <= 32'b11111100111110111111010011110011;
REG[5719] <= 32'b00011000000000111111110011111111;
REG[5720] <= 32'b11111110111100100001110100000111;
REG[5721] <= 32'b00000000111011111111011011101111;
REG[5722] <= 32'b00001000000000000001001011111000;
REG[5723] <= 32'b11110010111111011111100011110101;
REG[5724] <= 32'b00001011111100111111000100001000;
REG[5725] <= 32'b11110100111110010001001000010101;
REG[5726] <= 32'b00000001000001010000011000000010;
REG[5727] <= 32'b11111100111110111111101000001111;
REG[5728] <= 32'b00011000000000011111001111111110;
REG[5729] <= 32'b11111011000011110001001000000110;
REG[5730] <= 32'b11110011111101001111010000001011;
REG[5731] <= 32'b00000100000000010000000011111010;
REG[5732] <= 32'b00001011111100001111000111101111;
REG[5733] <= 32'b11110111111110100000011011110010;
REG[5734] <= 32'b11111111111101111111101111110001;
REG[5735] <= 32'b11110100111110111111111111111110;
REG[5736] <= 32'b11111001111110101111000011111000;
REG[5737] <= 32'b11110110000000101111010111111101;
REG[5738] <= 32'b00000101111110011111101011111001;
REG[5739] <= 32'b11110011111111110001011111110101;
REG[5740] <= 32'b11111010111111011110101111110010;
REG[5741] <= 32'b00000101000101110001011000000100;
REG[5742] <= 32'b11110001111100111111111111111001;
REG[5743] <= 32'b00000111000000111111100111110101;
REG[5744] <= 32'b11110110111110010000100111110011;
REG[5745] <= 32'b00000100000010110001000011110001;
REG[5746] <= 32'b11111110111100110000000111111111;
REG[5747] <= 32'b00000010111101100000101011110101;
REG[5748] <= 32'b11111011111100011111110011101110;
REG[5749] <= 32'b11110110111101001111100011111010;
REG[5750] <= 32'b11111010000000011111111100000010;
REG[5751] <= 32'b11111000111110111111001000000010;
REG[5752] <= 32'b11111011000001000000110100000111;
REG[5753] <= 32'b11110100000110010000100100001100;
REG[5754] <= 32'b00001101000100110001100011110110;
REG[5755] <= 32'b00000000111101100000010100010001;
REG[5756] <= 32'b00010100000001100000011011110101;
REG[5757] <= 32'b11111101111111000000000011111000;
REG[5758] <= 32'b11110110111101001111110100011011;
REG[5759] <= 32'b00010110111111011111101011100111;
REG[5760] <= 32'b11110110000111000000111100000111;
REG[5761] <= 32'b11111100111101010000001111111100;
REG[5762] <= 32'b11111000111111010000001100000000;
REG[5763] <= 32'b00000111111100111111100100001011;
REG[5764] <= 32'b00001100111111101111101111100110;
REG[5765] <= 32'b11101110000000000000100011111111;
REG[5766] <= 32'b00000101111011101110111100001101;
REG[5767] <= 32'b00001010000001011111111011101111;
REG[5768] <= 32'b11100101000001110000001000000010;
REG[5769] <= 32'b00000111111110101111000111110110;
REG[5770] <= 32'b00000011000010001111111111111010;
REG[5771] <= 32'b11111010111110101111111111111110;
REG[5772] <= 32'b00001001111101001111011011111011;
REG[5773] <= 32'b00001110000000001111110011101110;
REG[5774] <= 32'b11110001111110010001000011111011;
REG[5775] <= 32'b11111011111011111111100100000111;
REG[5776] <= 32'b00011111000011010000001111111101;
REG[5777] <= 32'b11110111000001010000000000001111;
REG[5778] <= 32'b11110101111011011111000000000100;
REG[5779] <= 32'b00000000000011111111101000001000;
REG[5780] <= 32'b11110101111110010000000100010100;
REG[5781] <= 32'b00010000000001110000011011110110;
REG[5782] <= 32'b11111010111101000000011111111101;
REG[5783] <= 32'b11111101111110010000001011111101;
REG[5784] <= 32'b00000111111111101110111111111010;
REG[5785] <= 32'b11111110111101010001100000001010;
REG[5786] <= 32'b00000011001101000001001100000110;
REG[5787] <= 32'b00001101000000110000011000010010;
REG[5788] <= 32'b00001101111101010001010011111100;
REG[5789] <= 32'b11111101000001001111011111111001;
REG[5790] <= 32'b00000100111111001111111011111010;
REG[5791] <= 32'b00001001111101100000100011111110;
REG[5792] <= 32'b11111001111111000001011111111100;
REG[5793] <= 32'b00001000111110110000010011111010;
REG[5794] <= 32'b11111101111100101111110111111111;
REG[5795] <= 32'b00000010111101101111110000000101;
REG[5796] <= 32'b00000101000010001111101011110110;
REG[5797] <= 32'b00000011000000110000010100000000;
REG[5798] <= 32'b00000000000000100001001100001100;
REG[5799] <= 32'b00000110111101111111011011110001;
REG[5800] <= 32'b00010000000000000000000011111000;
REG[5801] <= 32'b11110010111110010000100100000011;
REG[5802] <= 32'b11111010111100011110100100000001;
REG[5803] <= 32'b00001010000010001111101111110110;
REG[5804] <= 32'b11110011000010101111111100001001;
REG[5805] <= 32'b00000100111110101111010100001101;
REG[5806] <= 32'b00000010000011000000001111111010;
REG[5807] <= 32'b11111001000100000000001100001010;
REG[5808] <= 32'b00000011000000000000100011110001;
REG[5809] <= 32'b11101100111111011111101011111110;
REG[5810] <= 32'b11111111111101001111010000000111;
REG[5811] <= 32'b11101111111101001111011011111000;
REG[5812] <= 32'b11111000111101110000001011111011;
REG[5813] <= 32'b11110110000001101111110011101011;
REG[5814] <= 32'b00000001111101001111010100000011;
REG[5815] <= 32'b11111100111101011111001111111000;
REG[5816] <= 32'b11111000000001011111011111101011;
REG[5817] <= 32'b11110110111101111110111011111010;
REG[5818] <= 32'b11110111111010001111110100111001;
REG[5819] <= 32'b00101100111110001110110111011111;
REG[5820] <= 32'b11111101001001110001001111111110;
REG[5821] <= 32'b11111101111110000001100111111100;
REG[5822] <= 32'b00000000000001010000011011110111;
REG[5823] <= 32'b00001100111101011110111100010001;
REG[5824] <= 32'b00000111111111111111100000010000;
REG[5825] <= 32'b11111110111110111111011011111001;
REG[5826] <= 32'b11111000111101101111111000000110;
REG[5827] <= 32'b00000001111111101111010011101011;
REG[5828] <= 32'b11111011000000010001011000000001;
REG[5829] <= 32'b11110001111101000000001000000001;
REG[5830] <= 32'b00010001111111010001010000010101;
REG[5831] <= 32'b00000001000000110000001000010110;
REG[5832] <= 32'b00010000000101000000001111111001;
REG[5833] <= 32'b11111111000100111111011111110010;
REG[5834] <= 32'b11110011111110110000011100010111;
REG[5835] <= 32'b11111110000010101111101100001000;
REG[5836] <= 32'b00000011111110110000000000000000;
REG[5837] <= 32'b11111010000000101111111011111000;
REG[5838] <= 32'b00001010000010001111100011111001;
REG[5839] <= 32'b11111011111110100000010011111101;
REG[5840] <= 32'b11111010000010110001010100001010;
REG[5841] <= 32'b11111100111101101111101000001001;
REG[5842] <= 32'b00010010000001001111100011110011;
REG[5843] <= 32'b11111000000100110001001100010000;
REG[5844] <= 32'b11111010000001100000001000000100;
REG[5845] <= 32'b11111100000000010000001100001000;
REG[5846] <= 32'b11110000111110001111011011111101;
REG[5847] <= 32'b00000000001001011110111100000101;
REG[5848] <= 32'b00000001111111000000100000010001;
REG[5849] <= 32'b11111111000011000000001100001010;
REG[5850] <= 32'b11111000000001111111011000000011;
REG[5851] <= 32'b11111100000100001110110011101011;
REG[5852] <= 32'b11110100111111001110111111101100;
REG[5853] <= 32'b11110110000100010000101111110111;
REG[5854] <= 32'b11111000111101101111010100000101;
REG[5855] <= 32'b00000011111110100000000011111001;
REG[5856] <= 32'b00001110111110010000001111111010;
REG[5857] <= 32'b11111000111110000000111011110111;
REG[5858] <= 32'b11110010000000111111111011111100;
REG[5859] <= 32'b00101010000110000000001111111101;
REG[5860] <= 32'b11110011111110101111010011111100;
REG[5861] <= 32'b00000010111100101111001011110000;
REG[5862] <= 32'b00000010000000011111101111111110;
REG[5863] <= 32'b00001011000011100000011011111000;
REG[5864] <= 32'b11111101111111000000101100011000;
REG[5865] <= 32'b00011000111100011111000011110001;
REG[5866] <= 32'b11111010000001111111110111111010;
REG[5867] <= 32'b11111000000001000000110011111010;
REG[5868] <= 32'b11111101111011011111111100001111;
REG[5869] <= 32'b00101101111110101111011111110011;
REG[5870] <= 32'b00010010000001000000101111111100;
REG[5871] <= 32'b11111101000001100000001100010011;
REG[5872] <= 32'b00011001000010001111111011111100;
REG[5873] <= 32'b00000000000100010001000100001000;
REG[5874] <= 32'b00000111000100000000010100001001;
REG[5875] <= 32'b00011001000010000000011000000000;
REG[5876] <= 32'b11111001000001000000001111110010;
REG[5877] <= 32'b00000110111110001111100111111100;
REG[5878] <= 32'b00001000111110100000000111111101;
REG[5879] <= 32'b00000110111110000000001000000001;
REG[5880] <= 32'b00000000000001001111101100000100;
REG[5881] <= 32'b11111101000000010000001111111011;
REG[5882] <= 32'b00000000000010100000000011111010;
REG[5883] <= 32'b00011000000000011110110000001001;
REG[5884] <= 32'b11110110111101100001010100011001;
REG[5885] <= 32'b11110011111110011111100011110110;
REG[5886] <= 32'b00001100000010101111010111111101;
REG[5887] <= 32'b00000010111100101111111111111011;
REG[5888] <= 32'b11110101111101111111110111111011;
REG[5889] <= 32'b11111111111111010001001111110110;
REG[5890] <= 32'b11111011111111110000100011111110;
REG[5891] <= 32'b00001101111110011111011111111110;
REG[5892] <= 32'b00010111111110101111101011111100;
REG[5893] <= 32'b11111010111110101111110011110110;
REG[5894] <= 32'b11111010000001000000111000000010;
REG[5895] <= 32'b11110110111111010000010011111000;
REG[5896] <= 32'b11111110111110011111001100001100;
REG[5897] <= 32'b00000101111110111111101111111100;
REG[5898] <= 32'b11111010111111110000010111111100;
REG[5899] <= 32'b11110011111101111110111111101100;
REG[5900] <= 32'b00000000111101001110111111111000;
REG[5901] <= 32'b11110010111100000000001111111010;
REG[5902] <= 32'b11110111111101100001011100001100;
REG[5903] <= 32'b00000010111110111111010111100111;
REG[5904] <= 32'b00000101000000001111101100011111;
REG[5905] <= 32'b00010001111110111110111111110100;
REG[5906] <= 32'b11111011000010100001001000000100;
REG[5907] <= 32'b11111010111111111111101000000111;
REG[5908] <= 32'b00001100000010011111100111110110;
REG[5909] <= 32'b11110111000001110000010100000100;
REG[5910] <= 32'b11110011111101111111010100000100;
REG[5911] <= 32'b00000011000001110000100011111001;
REG[5912] <= 32'b11111000111110101111111011110111;
REG[5913] <= 32'b00000010111101101111100111110101;
REG[5914] <= 32'b11111100000000000000110011111011;
REG[5915] <= 32'b00000011111101011111110000001110;
REG[5916] <= 32'b11111110111111010001000100000011;
REG[5917] <= 32'b00001100111110001111000111111001;
REG[5918] <= 32'b00001011000011100001101011111100;
REG[5919] <= 32'b11111000111111000000111100000100;
REG[5920] <= 32'b00000111111110010000110100000011;
REG[5921] <= 32'b00010010000010010000100100001010;
REG[5922] <= 32'b00000111111110110000100000000101;
REG[5923] <= 32'b00000110000000110000101011111010;
REG[5924] <= 32'b00010000111111101111101000000110;
REG[5925] <= 32'b11111010000000101111100100000000;
REG[5926] <= 32'b11111100111101001111001111110100;
REG[5927] <= 32'b11110101111111011111101111110000;
REG[5928] <= 32'b11111001111101000000110100000001;
REG[5929] <= 32'b00000001111101110001111000000000;
REG[5930] <= 32'b11110111000001000000011100011011;
REG[5931] <= 32'b00010000000010101111101100000010;
REG[5932] <= 32'b00010000001010001111010000000000;
REG[5933] <= 32'b11111111111111111111111000011101;
REG[5934] <= 32'b00000111000011000001010011111001;
REG[5935] <= 32'b11111000111111100000011100000001;
REG[5936] <= 32'b00000001111101110000000000000101;
REG[5937] <= 32'b00001000000001110000001111110101;
REG[5938] <= 32'b11111001000000011111100000000000;
REG[5939] <= 32'b00000001111111111111110000000000;
REG[5940] <= 32'b11110111111100001111001011111010;
REG[5941] <= 32'b00000011000010010000000100000111;
REG[5942] <= 32'b11111101111110110000010000000111;
REG[5943] <= 32'b00000110000011100000010011111000;
REG[5944] <= 32'b11111100000011100000010111111111;
REG[5945] <= 32'b00000011000001000000110100010001;
REG[5946] <= 32'b00001001111110000000001111111111;
REG[5947] <= 32'b00001100000001000001000100001010;
REG[5948] <= 32'b11111011111111000000000100000110;
REG[5949] <= 32'b00000111111111111111011011101101;
REG[5950] <= 32'b11101110111101110000011011111101;
REG[5951] <= 32'b00000101111110011111010111111100;
REG[5952] <= 32'b11111001111111100000100011111011;
REG[5953] <= 32'b11110101111110101110010111100111;
REG[5954] <= 32'b00001100111111011111101011111001;
REG[5955] <= 32'b11110100111010011111011100000000;
REG[5956] <= 32'b11111011111101000001001000001010;
REG[5957] <= 32'b00001110000001110001000000000011;
REG[5958] <= 32'b00010000000110110000101111111111;
REG[5959] <= 32'b00000111000000110000111000001100;
REG[5960] <= 32'b00000011111111100000101111111100;
REG[5961] <= 32'b00000011111111001111100100000110;
REG[5962] <= 32'b00000101000001000001001000001011;
REG[5963] <= 32'b00000011000010011111111000000100;
REG[5964] <= 32'b11111110111111000000000000000111;
REG[5965] <= 32'b11111110000000101111101011110111;
REG[5966] <= 32'b11110101111111001111100111101111;
REG[5967] <= 32'b00000011111101001111010000000110;
REG[5968] <= 32'b00000111111110101111011111111000;
REG[5969] <= 32'b11111011111111101111101011110110;
REG[5970] <= 32'b11111000111111001111010011111110;
REG[5971] <= 32'b11111111000001111111100111111110;
REG[5972] <= 32'b11111011111110100000000111110110;
REG[5973] <= 32'b11110110111111110000010111111110;
REG[5974] <= 32'b00000111000000101111111011111010;
REG[5975] <= 32'b11101010000001010000010100000010;
REG[5976] <= 32'b00001011000101011111110000001101;
REG[5977] <= 32'b00000001111111110010000100100111;
REG[5978] <= 32'b11101110000011100000000100000011;
REG[5979] <= 32'b00000010000010010000010100000001;
REG[5980] <= 32'b00000011111111010000100000001111;
REG[5981] <= 32'b00011100111111000000011011111111;
REG[5982] <= 32'b11111101000001000001001011110110;
REG[5983] <= 32'b00000111000000100000101111110101;
REG[5984] <= 32'b11110111111100100001001100010111;
REG[5985] <= 32'b00001111111100111110010111101100;
REG[5986] <= 32'b00010011000101010001000100000100;
REG[5987] <= 32'b00000101111100010000011100001111;
REG[5988] <= 32'b11101110111100100000010100001000;
REG[5989] <= 32'b00000110000001011110011011101111;
REG[5990] <= 32'b00001101000001110000011100001010;
REG[5991] <= 32'b11101100111011011111110100000111;
REG[5992] <= 32'b00001011111111110000000011110110;
REG[5993] <= 32'b11111101111110011111011100000000;
REG[5994] <= 32'b11111101111011111111010011110110;
REG[5995] <= 32'b11111110111111100000010111110101;
REG[5996] <= 32'b00000000000000001111111111111110;
REG[5997] <= 32'b11110111111110011111110100000011;
REG[5998] <= 32'b00010001111111110000100011111001;
REG[5999] <= 32'b11101011111110110000011000000001;
REG[6000] <= 32'b00000110111110001110111111111011;
REG[6001] <= 32'b11111110000001101111010100000010;
REG[6002] <= 32'b00000000111111101111100100000010;
REG[6003] <= 32'b11111101000011101111100011101010;
REG[6004] <= 32'b11110000111101101111101100000001;
REG[6005] <= 32'b11111011111010101110110011111011;
REG[6006] <= 32'b11111011000000010000000111101110;
REG[6007] <= 32'b11101010111101101111011111111111;
REG[6008] <= 32'b00000010111110101110111111110111;
REG[6009] <= 32'b11111001111111110000010000000100;
REG[6010] <= 32'b11111010111101001111010111110110;
REG[6011] <= 32'b00000100000011100001100100001011;
REG[6012] <= 32'b11110001000001010000111100001110;
REG[6013] <= 32'b00110101000111111111010111110010;
REG[6014] <= 32'b11101010111100110000011000010010;
REG[6015] <= 32'b00010000000011010001000011111101;
REG[6016] <= 32'b11111100000001100001001000000011;
REG[6017] <= 32'b00001000000010100000001000000010;
REG[6018] <= 32'b00010000000000100000010011111111;
REG[6019] <= 32'b11111110111111000000011000000100;
REG[6020] <= 32'b11110010000000110000000111111001;
REG[6021] <= 32'b00000100000001111110111100010100;
REG[6022] <= 32'b00001010000000110000000100000100;
REG[6023] <= 32'b11110001000100100000100100000000;
REG[6024] <= 32'b00000000000001000000010000000101;
REG[6025] <= 32'b11111000111100100000010011111101;
REG[6026] <= 32'b11111011111111101110110011101010;
REG[6027] <= 32'b00000011111100101111000111111101;
REG[6028] <= 32'b11110011111100111111001111110011;
REG[6029] <= 32'b00000000111100100000001011111100;
REG[6030] <= 32'b11111101000000110000000011110000;
REG[6031] <= 32'b00001011000000000000001100000000;
REG[6032] <= 32'b00000011111110100000110111111110;
REG[6033] <= 32'b00001011000100000000001111111011;
REG[6034] <= 32'b00001000111111000000001111110010;
REG[6035] <= 32'b11110000111100101111010111111111;
REG[6036] <= 32'b11111001111001111111010000000001;
REG[6037] <= 32'b00000010111111110000010000000000;
REG[6038] <= 32'b00001000111111000000000000000011;
REG[6039] <= 32'b11111111111100000000000111110101;
REG[6040] <= 32'b11111110111111101111111011101111;
REG[6041] <= 32'b00000101111101101111111000000100;
REG[6042] <= 32'b00000100111110101111110100000010;
REG[6043] <= 32'b11111111111110100000000011111100;
REG[6044] <= 32'b11111101111111011111100111111010;
REG[6045] <= 32'b00000110000010010000010111110010;
REG[6046] <= 32'b11110011111110000000001000000101;
REG[6047] <= 32'b11111111111111010000011100001111;
REG[6048] <= 32'b00000001000000011111100011101100;
REG[6049] <= 32'b11110100111110111111110000000100;
REG[6050] <= 32'b11111100111110001111111000000010;
REG[6051] <= 32'b00000000000001110000010000001110;
REG[6052] <= 32'b11110000111111110000001111111110;
REG[6053] <= 32'b00000011000011010000110111111101;
REG[6054] <= 32'b00000001111110010000000011110100;
REG[6055] <= 32'b00000010000011100000000000000001;
REG[6056] <= 32'b11110111111110111111101011111100;
REG[6057] <= 32'b11110110111100101110100011111101;
REG[6058] <= 32'b11111010111110100000110000001001;
REG[6059] <= 32'b11111000000011101111111000000001;
REG[6060] <= 32'b11110111000000011111111100000101;
REG[6061] <= 32'b00001000111100011111010011110110;
REG[6062] <= 32'b11110110111110000000001011111111;
REG[6063] <= 32'b11101110111101001111111111110111;
REG[6064] <= 32'b11111110000000111111101011110000;
REG[6065] <= 32'b00000000000001010000101100000001;
REG[6066] <= 32'b11111001111011111111111011110101;
REG[6067] <= 32'b00001000000000111111010111110011;
REG[6068] <= 32'b00000011111101010000011000001100;
REG[6069] <= 32'b11111100111110100000001000000101;
REG[6070] <= 32'b11110101111110101111111100000000;
REG[6071] <= 32'b00000111000010000000011111111000;
REG[6072] <= 32'b11111001111111101111111111111101;
REG[6073] <= 32'b00000101111110101111100111111011;
REG[6074] <= 32'b11111000111111101111100111111010;
REG[6075] <= 32'b11111001111100111111011100000000;
REG[6076] <= 32'b11111111111111011111110111110000;
REG[6077] <= 32'b11111001111110010000000111111101;
REG[6078] <= 32'b00000101000010111111101100000001;
REG[6079] <= 32'b00000000111110111111110011110001;
REG[6080] <= 32'b11110100000000001111100111110011;
REG[6081] <= 32'b11110001111011011110111100000110;
REG[6082] <= 32'b11111100000011100000001000010100;
REG[6083] <= 32'b11100010000010000001011100010001;
REG[6084] <= 32'b00000101001001111110111000001001;
REG[6085] <= 32'b00011010000110111110100000001100;
REG[6086] <= 32'b11101001000001110010011100100110;
REG[6087] <= 32'b11111100111111101111011111110110;
REG[6088] <= 32'b00000010000000001111111111111110;
REG[6089] <= 32'b11110110111101101111100011111000;
REG[6090] <= 32'b00000101111111011111111111111111;
REG[6091] <= 32'b11111100111110100001101000001101;
REG[6092] <= 32'b00000010000000100000001000001010;
REG[6093] <= 32'b00010111001001010001000100010110;
REG[6094] <= 32'b00100000000101100001011000011000;
REG[6095] <= 32'b00001100000010110001110100010111;
REG[6096] <= 32'b00000100111111110001001011110011;
REG[6097] <= 32'b11111100111110010000101000001000;
REG[6098] <= 32'b00001000111010111111111011101110;
REG[6099] <= 32'b00000011111111101111000111101111;
REG[6100] <= 32'b00000101111100011111101011111001;
REG[6101] <= 32'b11110001000101010001101000000001;
REG[6102] <= 32'b00000000111110001111011000000010;
REG[6103] <= 32'b00010010000011111111011011110000;
REG[6104] <= 32'b11110100000000010000000011110100;
REG[6105] <= 32'b00010010111100111111011111101110;
REG[6106] <= 32'b11110001111111000001010011101110;
REG[6107] <= 32'b11110100000010100000110000000111;
REG[6108] <= 32'b00001010111100011111100011111001;
REG[6109] <= 32'b11111110000011001111011111111011;
REG[6110] <= 32'b00010000111111110000100100000111;
REG[6111] <= 32'b11110011111101110000011100000101;
REG[6112] <= 32'b00010010000011110000100111111101;
REG[6113] <= 32'b00001011000101010001000100000011;
REG[6114] <= 32'b11111101000001000000001100000000;
REG[6115] <= 32'b00000010111111111111110100001000;
REG[6116] <= 32'b00001001000001011111101011111100;
REG[6117] <= 32'b11110110111111010000100000000000;
REG[6118] <= 32'b11111011111110111111100111111011;
REG[6119] <= 32'b00000000111111101111101011111010;
REG[6120] <= 32'b00000000000110011111111100000100;
REG[6121] <= 32'b00001101000101001111001000000111;
REG[6122] <= 32'b11110010111111010000001100001000;
REG[6123] <= 32'b00001100111111100000011011111110;
REG[6124] <= 32'b11111010111011000001000000000000;
REG[6125] <= 32'b11110111000001000000101100000011;
REG[6126] <= 32'b00000101111110001110011100001000;
REG[6127] <= 32'b00001001000001011111011011110101;
REG[6128] <= 32'b11110010111011010000100100010011;
REG[6129] <= 32'b11111011111101011111000111110010;
REG[6130] <= 32'b00000110000011111111101111110100;
REG[6131] <= 32'b11110101111101000000000000001100;
REG[6132] <= 32'b11111100000010110000101100000010;
REG[6133] <= 32'b11110101111110100000010100001001;
REG[6134] <= 32'b00000100000000011111101111111011;
REG[6135] <= 32'b00001011000001000000001100000010;
REG[6136] <= 32'b00000110111101010000000000000000;
REG[6137] <= 32'b00000101000010100000100000000011;
REG[6138] <= 32'b11111100000001010000011111111101;
REG[6139] <= 32'b00000100111111110000000111111100;
REG[6140] <= 32'b11110110111011111111001111110001;
REG[6141] <= 32'b00000011000000001110110100001011;
REG[6142] <= 32'b00010010000000110000100000001011;
REG[6143] <= 32'b11101010111111001111111111111000;
REG[6144] <= 32'b00010010000100011111011111111010;
REG[6145] <= 32'b11111001111110011111100011111011;
REG[6146] <= 32'b11111110111110001111010111111000;
REG[6147] <= 32'b11111010111111011111001111111100;
REG[6148] <= 32'b11110010111110001111111111111000;
REG[6149] <= 32'b11110010000011100000100011111100;
REG[6150] <= 32'b00000010111110010000011011101011;
REG[6151] <= 32'b00000000000010000000001111111110;
REG[6152] <= 32'b11110001111011110001001100001111;
REG[6153] <= 32'b11111011000001111111001011110010;
REG[6154] <= 32'b11110100000000100000000100001001;
REG[6155] <= 32'b00011100111101101111101111110111;
REG[6156] <= 32'b00000100000001110001110011111001;
REG[6157] <= 32'b11111110111100011111101100001000;
REG[6158] <= 32'b00001111000000000000000111111110;
REG[6159] <= 32'b00000101000000001111011000000110;
REG[6160] <= 32'b11111111000101110001000100001011;
REG[6161] <= 32'b11111010000001001111100000001011;
REG[6162] <= 32'b00001010000100000000000100001010;
REG[6163] <= 32'b00000101000101000001011000010110;
REG[6164] <= 32'b00000111111110110000100111111110;
REG[6165] <= 32'b00001000000000101111100011110010;
REG[6166] <= 32'b00000011111111100010010000010100;
REG[6167] <= 32'b00001001111111110000100000000001;
REG[6168] <= 32'b11111110111101011111100011110010;
REG[6169] <= 32'b11101010111101000001000011110111;
REG[6170] <= 32'b11110110111011101111001011110011;
REG[6171] <= 32'b00011100000010001111011011110010;
REG[6172] <= 32'b00000110000000101111110111110111;
REG[6173] <= 32'b11111000111100000000000011111110;
REG[6174] <= 32'b11110010111100011110110011101010;
REG[6175] <= 32'b11110001111101101110111111111000;
REG[6176] <= 32'b11111001111101101111111011111011;
REG[6177] <= 32'b00000000000000011111111111110110;
REG[6178] <= 32'b00000110000010001111111111111000;
REG[6179] <= 32'b11110101111100111111110000000010;
REG[6180] <= 32'b11111010111101110000000111111011;
REG[6181] <= 32'b11111111000000111111010011110100;
REG[6182] <= 32'b00000001111111111111101111111001;
REG[6183] <= 32'b11110000111110011111110111110111;
REG[6184] <= 32'b11110110111101111111001011111100;
REG[6185] <= 32'b00000011111101001110111111110010;
REG[6186] <= 32'b00001100000110000000000100000011;
REG[6187] <= 32'b00001100000000110000111000001001;
REG[6188] <= 32'b11111100000000110000010100000001;
REG[6189] <= 32'b00001010111111101111001000000010;
REG[6190] <= 32'b00000111111111001111001011101111;
REG[6191] <= 32'b11110011111100101111001011110001;
REG[6192] <= 32'b11110011111011011110111011111001;
REG[6193] <= 32'b11111101111101101111101111111101;
REG[6194] <= 32'b11111010000000011111110111111011;
REG[6195] <= 32'b00000111111111100001001000000111;
REG[6196] <= 32'b11110011111111000000001100000000;
REG[6197] <= 32'b00001100000011011111111011111111;
REG[6198] <= 32'b11111000111101001111111100001110;
REG[6199] <= 32'b00000001111111100001000100000000;
REG[6200] <= 32'b11110110000001111111110111110100;
REG[6201] <= 32'b00001111000000001111010100000101;
REG[6202] <= 32'b11111110111101000000111011111001;
REG[6203] <= 32'b11101101111111011111111111111100;
REG[6204] <= 32'b00001111000011011111011011110111;
REG[6205] <= 32'b11111001111101000000011100010111;
REG[6206] <= 32'b00000000111010001111111011110000;
REG[6207] <= 32'b11111101000010110000010011101100;
REG[6208] <= 32'b11110110111111010000011111110011;
REG[6209] <= 32'b00000011000001001111111100000000;
REG[6210] <= 32'b00000111111111100000100000000101;
REG[6211] <= 32'b11111111111111000000000000000011;
REG[6212] <= 32'b00001001000010111111110011111100;
REG[6213] <= 32'b00000111111011111111000100000001;
REG[6214] <= 32'b11111010000000100000101011110011;
REG[6215] <= 32'b11110001000000101111101000000001;
REG[6216] <= 32'b00011100000000001110011111110110;
REG[6217] <= 32'b11111110111111000000001000000100;
REG[6218] <= 32'b00001110111100111111111000000011;
REG[6219] <= 32'b11111011111110100001000011110000;
REG[6220] <= 32'b11111111000001010000001100000101;
REG[6221] <= 32'b00001001111100101111110000000011;
REG[6222] <= 32'b11110001111101100010010000000110;
REG[6223] <= 32'b00000111111110111111000011101011;
REG[6224] <= 32'b00000000000000101111111111110100;
REG[6225] <= 32'b11110001111100000000010111111111;
REG[6226] <= 32'b00000101111110001110110100000011;
REG[6227] <= 32'b11111011000010010001000000001011;
REG[6228] <= 32'b11110011000111111111110011111101;
REG[6229] <= 32'b11111000111111001111000000011000;
REG[6230] <= 32'b00000001000011000000001111101110;
REG[6231] <= 32'b11111011111101001111100100000011;
REG[6232] <= 32'b11111010111111111111110011111010;
REG[6233] <= 32'b11101110111011001110111111111001;
REG[6234] <= 32'b11110010111101101111010011110111;
REG[6235] <= 32'b00000000000011111111010000001001;
REG[6236] <= 32'b11110100111111001111100100000000;
REG[6237] <= 32'b00000010000101110000000011111111;
REG[6238] <= 32'b00000010000001001111100100001110;
REG[6239] <= 32'b11111001000010110001011000010010;
REG[6240] <= 32'b11110001111010101110111100001010;
REG[6241] <= 32'b11111001111111111110101111100100;
REG[6242] <= 32'b11110010000100011111111100000110;
REG[6243] <= 32'b11110101111011011111101000010100;
REG[6244] <= 32'b00000000000010010001001100001110;
REG[6245] <= 32'b00000111111110100000010111111101;
REG[6246] <= 32'b00010101000100010000010000000010;
REG[6247] <= 32'b00000010111111110001000100000010;
REG[6248] <= 32'b11111111111110011111101111111001;
REG[6249] <= 32'b00001110000010110000001111111110;
REG[6250] <= 32'b11110111111100000000100000000011;
REG[6251] <= 32'b11110111000001011111011011101001;
REG[6252] <= 32'b11110110111110011111110011111101;
REG[6253] <= 32'b11110000111010000001000111111111;
REG[6254] <= 32'b00001001000100010000010111101001;
REG[6255] <= 32'b00000010111101001111100111100100;
REG[6256] <= 32'b11101101111111001111000111111011;
REG[6257] <= 32'b11111000111110100000111100011100;
REG[6258] <= 32'b00010001000001101111101011101100;
REG[6259] <= 32'b11111011111100001111111000000100;
REG[6260] <= 32'b11111111000010010000101111110111;
REG[6261] <= 32'b11110101111111111111110100001100;
REG[6262] <= 32'b00001010111101010000011000000111;
REG[6263] <= 32'b00001010111101011111000111110100;
REG[6264] <= 32'b11111110000000101111101111110111;
REG[6265] <= 32'b11110101111110010000110100001011;
REG[6266] <= 32'b00000100111111101111010000000110;
REG[6267] <= 32'b00000000111110110000000000000010;
REG[6268] <= 32'b00000100111101001111111111111100;
REG[6269] <= 32'b00000001000010010001010000000000;
REG[6270] <= 32'b11111010111101011111011011111111;
REG[6271] <= 32'b11111111111100110000000000000111;
REG[6272] <= 32'b00000010111101101111100000001110;
REG[6273] <= 32'b00001110000001011111011011111100;
REG[6274] <= 32'b11110111000001100000100000010001;
REG[6275] <= 32'b00001001000000010000010100000110;
REG[6276] <= 32'b00000000111110011111010111111001;
REG[6277] <= 32'b11100100000011110000011000000010;
REG[6278] <= 32'b00000000000000101110101100001101;
REG[6279] <= 32'b00010000000001000000001011111100;
REG[6280] <= 32'b11101011000011100001011100100101;
REG[6281] <= 32'b11111011000000011111111111110110;
REG[6282] <= 32'b11110111000001111111011011110111;
REG[6283] <= 32'b11101001000001011111011111101100;
REG[6284] <= 32'b00000001000010100000100000000001;
REG[6285] <= 32'b11111000111110010000000111110110;
REG[6286] <= 32'b11111110111101111111110011110101;
REG[6287] <= 32'b00000001000000100000111111110111;
REG[6288] <= 32'b00001000111110110000011000001011;
REG[6289] <= 32'b00010001111111000000011100010101;
REG[6290] <= 32'b00010100000000111111111111111100;
REG[6291] <= 32'b00010011000011100000010100000001;
REG[6292] <= 32'b11110101111110000000100111111110;
REG[6293] <= 32'b00001010000110001111111111101111;
REG[6294] <= 32'b00001111000001101111011011111110;
REG[6295] <= 32'b00000000111011101111100011111111;
REG[6296] <= 32'b11110000000010000001001111111011;
REG[6297] <= 32'b11111011000000011111011011111011;
REG[6298] <= 32'b00000101111111100000000111101111;
REG[6299] <= 32'b11111011111101101111001111101101;
REG[6300] <= 32'b00001100111111011111010000000100;
REG[6301] <= 32'b00000111111100010000011011111110;
REG[6302] <= 32'b11110101000011110000111111111100;
REG[6303] <= 32'b00001001000100100000010011110010;
REG[6304] <= 32'b11111111111101110000011000010010;
REG[6305] <= 32'b11111111111110110000001111111111;
REG[6306] <= 32'b11111100000001011111101111111010;
REG[6307] <= 32'b00000100000000001110111111111001;
REG[6308] <= 32'b11111011000000000000000000000001;
REG[6309] <= 32'b11110100111110001111110100000001;
REG[6310] <= 32'b00000001000001011111000111110011;
REG[6311] <= 32'b11110111000011100000110000000001;
REG[6312] <= 32'b00010110000011101110011011111110;
REG[6313] <= 32'b11111001000001100010000100100001;
REG[6314] <= 32'b11110111111111110000101100000101;
REG[6315] <= 32'b00001001000010011111000000001011;
REG[6316] <= 32'b00001000000001010001111000001100;
REG[6317] <= 32'b11110111111101111111101100001101;
REG[6318] <= 32'b00001110111110001111011111110011;
REG[6319] <= 32'b11110110000010100000100100001110;
REG[6320] <= 32'b00000001000000001111110000001011;
REG[6321] <= 32'b11111101111101110000011000000000;
REG[6322] <= 32'b11111101000001011111111111111000;
REG[6323] <= 32'b00000101000010101111111111111110;
REG[6324] <= 32'b00001000111111010000011100001000;
REG[6325] <= 32'b00000010111111100000101000000100;
REG[6326] <= 32'b11111001111100110000000111110001;
REG[6327] <= 32'b00001110111110111111110000000100;
REG[6328] <= 32'b00000010000001110001011000000111;
REG[6329] <= 32'b00001000000101100000111000000110;
REG[6330] <= 32'b11111101111111111111101111111110;
REG[6331] <= 32'b11101010111011011111101011111101;
REG[6332] <= 32'b11111100000000101111001011101100;
REG[6333] <= 32'b00000000000001010000001100000011;
REG[6334] <= 32'b11111000111101110000001100000010;
REG[6335] <= 32'b11111001000110100000000111110100;
REG[6336] <= 32'b00000010000001100000011000010100;
REG[6337] <= 32'b00000110111110101111110000000101;
REG[6338] <= 32'b00001110000000110000010000000010;
REG[6339] <= 32'b11110100111101110000011111101110;
REG[6340] <= 32'b00001001111111101111011011111111;
REG[6341] <= 32'b00001000111110100000111100001001;
REG[6342] <= 32'b11111001111110000000001011101110;
REG[6343] <= 32'b11110111000000101111001011111000;
REG[6344] <= 32'b11110010111010101111101100000000;
REG[6345] <= 32'b00000000111111100000001111110010;
REG[6346] <= 32'b11111010111110001111101000000011;
REG[6347] <= 32'b00000011111101101111110011111110;
REG[6348] <= 32'b00000010000101110000000111110000;
REG[6349] <= 32'b00010110111010110000010100011110;
REG[6350] <= 32'b00000011111011000000101011101010;
REG[6351] <= 32'b11111010000010001111110011100111;
REG[6352] <= 32'b00000110111011011111110000000110;
REG[6353] <= 32'b00001100111110001111111100000000;
REG[6354] <= 32'b11110100000000000000000011110101;
REG[6355] <= 32'b11110100111111000000000111111101;
REG[6356] <= 32'b00000100111101111111101000000010;
REG[6357] <= 32'b00001001000001100000101011101110;
REG[6358] <= 32'b11110011111110000000101000000011;
REG[6359] <= 32'b11111110111110000000000111110001;
REG[6360] <= 32'b00001001000001110000000011111110;
REG[6361] <= 32'b11111110111101000001010000000011;
REG[6362] <= 32'b11110110000100010000110000000001;
REG[6363] <= 32'b00010110111100101111001011111101;
REG[6364] <= 32'b00000111111111010001000011110111;
REG[6365] <= 32'b11110011111110000000011100010110;
REG[6366] <= 32'b00000001000110000001001000000101;
REG[6367] <= 32'b11111000111100101111001000001001;
REG[6368] <= 32'b00000110000010010000011111111010;
REG[6369] <= 32'b11111101111111100000001000000011;
REG[6370] <= 32'b00000100111111011111110011110001;
REG[6371] <= 32'b11110110111110001111010011101110;
REG[6372] <= 32'b11111100111101001111100111111011;
REG[6373] <= 32'b11111110111100000000000000000000;
REG[6374] <= 32'b00000100000100001111110111110000;
REG[6375] <= 32'b00010100000110100000001011101100;
REG[6376] <= 32'b11110100111001100000100000001100;
REG[6377] <= 32'b11111001000000010000000111111001;
REG[6378] <= 32'b11111100000001100000001100010010;
REG[6379] <= 32'b00001010111111010000110100001010;
REG[6380] <= 32'b00001100111110111111001011101100;
REG[6381] <= 32'b00000100000010110000100100000110;
REG[6382] <= 32'b11110010111101011111010011111101;
REG[6383] <= 32'b11111010000000001111010111110101;
REG[6384] <= 32'b00000100000000011111101111111110;
REG[6385] <= 32'b11110111000010100000111000001011;
REG[6386] <= 32'b11111101111111110000001000000010;
REG[6387] <= 32'b00100000000010111111100100010000;
REG[6388] <= 32'b00001011000000000000010100000010;
REG[6389] <= 32'b11110010111101010000010011110101;
REG[6390] <= 32'b11110010000001111111111011110000;
REG[6391] <= 32'b00000000000001101111101000000111;
REG[6392] <= 32'b00000011111011011111001111111010;
REG[6393] <= 32'b11110101000001001111110100011011;
REG[6394] <= 32'b11101011111101110000000111111001;
REG[6395] <= 32'b11110100000101111111000011110100;
REG[6396] <= 32'b00000001000000010000001100000000;
REG[6397] <= 32'b00000110111111001111010000000010;
REG[6398] <= 32'b00001100111101111111110111101011;
REG[6399] <= 32'b11110011111101100000001100010111;
REG[6400] <= 32'b00011101000000101111001111111010;
REG[6401] <= 32'b00001001111101011110111011101111;
REG[6402] <= 32'b00000100000000000000010000001100;
REG[6403] <= 32'b00000000000011111111110011111010;
REG[6404] <= 32'b11111001000010111111011111110110;
REG[6405] <= 32'b11110111111110000000010100000010;
REG[6406] <= 32'b00000100111110110000010000000011;
REG[6407] <= 32'b00000000111111100000000100000101;
REG[6408] <= 32'b00001000111101000000110000000010;
REG[6409] <= 32'b11110111000000010000010011110100;
REG[6410] <= 32'b00001100111110101111010000000100;
REG[6411] <= 32'b11111101000011010000001111111001;
REG[6412] <= 32'b11111001000010100010000100110110;
REG[6413] <= 32'b00101000111111000000000011110110;
REG[6414] <= 32'b00001110000100110000101011110111;
REG[6415] <= 32'b11111011111011101111100111110111;
REG[6416] <= 32'b00001010000001111111110011111101;
REG[6417] <= 32'b11111000111111000000011100000000;
REG[6418] <= 32'b00001000000010101111111011111110;
REG[6419] <= 32'b00000000111110000000111100000001;
REG[6420] <= 32'b11100111111100001111111011111000;
REG[6421] <= 32'b11101010000110100000011100000010;
REG[6422] <= 32'b11110101111101011110100000000011;
REG[6423] <= 32'b11110101111110001110001111111010;
REG[6424] <= 32'b11101110000000011111010111101110;
REG[6425] <= 32'b11110100111110001111000111111011;
REG[6426] <= 32'b00000111000000001111101011110011;
REG[6427] <= 32'b00000100001001100000010011111100;
REG[6428] <= 32'b00000001000000100000010000001010;
REG[6429] <= 32'b00001001000100010001001100001001;
REG[6430] <= 32'b00010000000011010000000111111010;
REG[6431] <= 32'b11110011000101000010001100000101;
REG[6432] <= 32'b00000110000000111111001111111100;
REG[6433] <= 32'b11110111111100111111100011110110;
REG[6434] <= 32'b11110000111111100000011100000000;
REG[6435] <= 32'b11101011111101011111000000010110;
REG[6436] <= 32'b00000110000001011111000111110111;
REG[6437] <= 32'b11101111000011001111111100010010;
REG[6438] <= 32'b11111010111101101111001011110111;
REG[6439] <= 32'b00000101000010011111100111111001;
REG[6440] <= 32'b11101101000000010000100011111101;
REG[6441] <= 32'b11111010111101111110110100000101;
REG[6442] <= 32'b00000101111111101111001011111110;
REG[6443] <= 32'b00000101000001010000110111111110;
REG[6444] <= 32'b11101100000001100001001100001011;
REG[6445] <= 32'b00010000000000101111010000000011;
REG[6446] <= 32'b00001101000000100001000100001110;
REG[6447] <= 32'b11111101000000101111111011110010;
REG[6448] <= 32'b11110100111110001110111100001000;
REG[6449] <= 32'b00001100111100001110101111110000;
REG[6450] <= 32'b11101111111110111111110011111010;
REG[6451] <= 32'b11110110111011001111001000000010;
REG[6452] <= 32'b00001100000000101111000011110110;
REG[6453] <= 32'b11101110111111110000111000000010;
REG[6454] <= 32'b11101110111101101111000111111111;
REG[6455] <= 32'b00001010000001111111000111111001;
REG[6456] <= 32'b00000111000010010001010011111111;
REG[6457] <= 32'b11101111111100101111111011111000;
REG[6458] <= 32'b00001010000001100010101000001101;
REG[6459] <= 32'b11111011111011101110110011110011;
REG[6460] <= 32'b11110000000001111111001011110001;
REG[6461] <= 32'b11111111111100001110001111111110;
REG[6462] <= 32'b11101101111101000000110011110010;
REG[6463] <= 32'b00001011001100011111000111110010;
REG[6464] <= 32'b00000101111010111111101000010101;
REG[6465] <= 32'b11110110111101111111011100010110;
REG[6466] <= 32'b00000110000000001111110111110100;
REG[6467] <= 32'b11110110000010101111101100000001;
REG[6468] <= 32'b00010100000010001111000100010001;
REG[6469] <= 32'b00000111000100001111100000000000;
REG[6470] <= 32'b00000000000000100000000000001101;
REG[6471] <= 32'b11111011111111001111010011111101;
REG[6472] <= 32'b11111001000001001111010111110110;
REG[6473] <= 32'b11110111111110011111000111110111;
REG[6474] <= 32'b11111111111110100000010000001101;
REG[6475] <= 32'b00001010000100101111111000000000;
REG[6476] <= 32'b00000000111111001111010100001101;
REG[6477] <= 32'b00000100111100111110100111110111;
REG[6478] <= 32'b11111000000000101111101111110111;
REG[6479] <= 32'b11111110111100101111010111101011;
REG[6480] <= 32'b11110111111110010000000000001011;
REG[6481] <= 32'b00000101111111111111101011111011;
REG[6482] <= 32'b00000001000010110000100000000100;
REG[6483] <= 32'b00000011000000000000101011111100;
REG[6484] <= 32'b00000001111101011111001111111000;
REG[6485] <= 32'b11111111000001101111111111111011;
REG[6486] <= 32'b11110000111111000000000111111101;
REG[6487] <= 32'b11110110111110111111100111111101;
REG[6488] <= 32'b00000001000001011111011100000001;
REG[6489] <= 32'b11110100111101011111100100001001;
REG[6490] <= 32'b11111100111101111111010011111110;
REG[6491] <= 32'b11111101111110001111011111110101;
REG[6492] <= 32'b00001111111111111111001111100101;
REG[6493] <= 32'b11111101111111110000100100000010;
REG[6494] <= 32'b00000011111100111111111011111101;
REG[6495] <= 32'b00001000111110101111100000001000;
REG[6496] <= 32'b00000101111111111111111011111111;
REG[6497] <= 32'b00000001000000101111001111110111;
REG[6498] <= 32'b11111101000110000000011111110101;
REG[6499] <= 32'b11101110111110001111011100001011;
REG[6500] <= 32'b00000101111100001110101111110001;
REG[6501] <= 32'b11111100111111001111111100000001;
REG[6502] <= 32'b11110100111110011110101011110000;
REG[6503] <= 32'b00001010111011101111001111110011;
REG[6504] <= 32'b11111100111011100000010111111001;
REG[6505] <= 32'b11111010111100110000001111111110;
REG[6506] <= 32'b00000111000000010000000111110000;
REG[6507] <= 32'b11111101111111110000001100000001;
REG[6508] <= 32'b00010000000011000000001000000100;
REG[6509] <= 32'b00000100111111110000111100001010;
REG[6510] <= 32'b11111101111101011110110000000101;
REG[6511] <= 32'b00000100000100011111011011110010;
REG[6512] <= 32'b11111010000001000000001100001011;
REG[6513] <= 32'b11111100111100110000001000001010;
REG[6514] <= 32'b00010110000101001111110000000011;
REG[6515] <= 32'b00000001111101101111101111111010;
REG[6516] <= 32'b11111101000010010001011111101111;
REG[6517] <= 32'b11111111111110111111100000001001;
REG[6518] <= 32'b00001101111100000000000111111011;
REG[6519] <= 32'b00010110111111100000010100000111;
REG[6520] <= 32'b00001010111111011111110111110100;
REG[6521] <= 32'b11111100000011100000010000000010;
REG[6522] <= 32'b11110000111101101111010100010110;
REG[6523] <= 32'b00000111000010000000010000000101;
REG[6524] <= 32'b00001000000100101111010111111010;
REG[6525] <= 32'b11110101111111100000110100001110;
REG[6526] <= 32'b11110001111110011111111011111010;
REG[6527] <= 32'b00001100000101111111100000000001;
REG[6528] <= 32'b00000101000001011111111000010101;
REG[6529] <= 32'b00001000000000111111101100000000;
REG[6530] <= 32'b11111011000011100001001100001001;
REG[6531] <= 32'b11110101111110111111011111110111;
REG[6532] <= 32'b00001110111111111111111111111101;
REG[6533] <= 32'b11111101111010011111100011111001;
REG[6534] <= 32'b00001111000000100001110111100111;
REG[6535] <= 32'b11101100111101100000010000000000;
REG[6536] <= 32'b00011111111100101111000011111011;
REG[6537] <= 32'b11111001000010100000011111111001;
REG[6538] <= 32'b11101110000000111111110111110001;
REG[6539] <= 32'b11100100000000101111101111110100;
REG[6540] <= 32'b11111011000000011111111000010101;
REG[6541] <= 32'b00001000111110101111101111110110;
REG[6542] <= 32'b11101011000010011111001111110000;
REG[6543] <= 32'b00000111111111010001001000001100;
REG[6544] <= 32'b11110101111011000000010000001000;
REG[6545] <= 32'b00001101111101101111101111110011;
REG[6546] <= 32'b11111001111101101111011000000110;
REG[6547] <= 32'b11111001111010100000110011111011;
REG[6548] <= 32'b11101110000010111111010111111001;
REG[6549] <= 32'b00000010111111011111000111111110;
REG[6550] <= 32'b11111010000000010000001100000011;
REG[6551] <= 32'b00000110111010110000101011110110;
REG[6552] <= 32'b00000001111101001111000000000011;
REG[6553] <= 32'b00101011111111010000011011110110;
REG[6554] <= 32'b11101000111101100000101111101001;
REG[6555] <= 32'b11110101111110101111111100001110;
REG[6556] <= 32'b00100111000101011111011011110000;
REG[6557] <= 32'b11111100000100100001110000101000;
REG[6558] <= 32'b11111110111111010000011011111111;
REG[6559] <= 32'b11111101111110110000111111111110;
REG[6560] <= 32'b11111010000011100000010100000010;
REG[6561] <= 32'b11111110000000000001110000010111;
REG[6562] <= 32'b00010010000010001111100000000110;
REG[6563] <= 32'b00011010000010000000010000000011;
REG[6564] <= 32'b00000000000010000001001000001100;
REG[6565] <= 32'b11101000111101011111100011110000;
REG[6566] <= 32'b00000001111101101111010100000000;
REG[6567] <= 32'b00000001000010100000111011111010;
REG[6568] <= 32'b00000000000010100000000111111010;
REG[6569] <= 32'b11110001111111110000000100001101;
REG[6570] <= 32'b00000100000000111111000000000000;
REG[6571] <= 32'b11111111000010110001010000000001;
REG[6572] <= 32'b11111101000000110000010100001000;
REG[6573] <= 32'b00000110000000110001001111110110;
REG[6574] <= 32'b11110110111011101111100011110011;
REG[6575] <= 32'b00000001000001101111110111110000;
REG[6576] <= 32'b11101111111010101111010100001000;
REG[6577] <= 32'b00010101000100111111101011110111;
REG[6578] <= 32'b11111000111111011111110011110100;
REG[6579] <= 32'b00000110111101001111110100001001;
REG[6580] <= 32'b00011111111101000000010111110111;
REG[6581] <= 32'b11101010111100110000111011111110;
REG[6582] <= 32'b00000101111100011111000111110100;
REG[6583] <= 32'b00010011000100011111111111111101;
REG[6584] <= 32'b11101111111101110001011100001111;
REG[6585] <= 32'b11111111111111101111011111111010;
REG[6586] <= 32'b00000110000011010000001000000100;
REG[6587] <= 32'b11111010111111001111011111110000;
REG[6588] <= 32'b00000101111111110000100111111101;
REG[6589] <= 32'b11110000111100001111101011110111;
REG[6590] <= 32'b11111100000010101111011011110110;
REG[6591] <= 32'b00001010111100001111011011101111;
REG[6592] <= 32'b11110100111101010000111111111001;
REG[6593] <= 32'b11111111111101101111111111111001;
REG[6594] <= 32'b00001110000001110000110111111010;
REG[6595] <= 32'b00001000000000111111111000000110;
REG[6596] <= 32'b11110110111101101110111000000010;
REG[6597] <= 32'b00000001111111011111100000000100;
REG[6598] <= 32'b00000000000001010000000000000000;
REG[6599] <= 32'b11111011000001011111100000001000;
REG[6600] <= 32'b00000010111111000000101111011000;
REG[6601] <= 32'b00010101111111110000000111110001;
REG[6602] <= 32'b11110101000011000001101011101111;
REG[6603] <= 32'b00000000111110001111110011111100;
REG[6604] <= 32'b11110011111010110000100100001111;
REG[6605] <= 32'b11110111111110100010011111111101;
REG[6606] <= 32'b11111100111110001110101111111111;
REG[6607] <= 32'b01000010000001110000001111111010;
REG[6608] <= 32'b11110011111110100001001011110000;
REG[6609] <= 32'b11111111000010110000110000001011;
REG[6610] <= 32'b00001111111110111111011111110011;
REG[6611] <= 32'b11111010111110110000001011110011;
REG[6612] <= 32'b00000101111111110000100011101101;
REG[6613] <= 32'b11110000111100101111101011110111;
REG[6614] <= 32'b11110011000000101111011000000110;
REG[6615] <= 32'b11111000111110011111001011111100;
REG[6616] <= 32'b11101011000000111111000111110011;
REG[6617] <= 32'b11110100000000111111001100000111;
REG[6618] <= 32'b11111110111101111111011011111100;
REG[6619] <= 32'b11111111111100011111010111110101;
REG[6620] <= 32'b11110100000001010000100111110011;
REG[6621] <= 32'b11111010111110011111100000000110;
REG[6622] <= 32'b00000101111111110000000011111011;
REG[6623] <= 32'b11101111111100101111110011111011;
REG[6624] <= 32'b00000101000001100000011100000000;
REG[6625] <= 32'b00000100000010000000111100000100;
REG[6626] <= 32'b00000000000000111111101000000000;
REG[6627] <= 32'b11111111111111110000101111111100;
REG[6628] <= 32'b00000001111110010000010111111100;
REG[6629] <= 32'b00001011111101110000001000000100;
REG[6630] <= 32'b11111000111101101111100100001010;
REG[6631] <= 32'b00000101111111111111011100000110;
REG[6632] <= 32'b00001111111101111110011111110001;
REG[6633] <= 32'b11111101000001001111111011111110;
REG[6634] <= 32'b11101100111101001111000111111100;
REG[6635] <= 32'b11101110111110011110110011110000;
REG[6636] <= 32'b00010001111110101111011111111010;
REG[6637] <= 32'b11110111000010000001000000010100;
REG[6638] <= 32'b11111010111110011111110100001111;
REG[6639] <= 32'b00000110000010010000001000000000;
REG[6640] <= 32'b00010001000001011111101011111101;
REG[6641] <= 32'b00001001111110001111110011111110;
REG[6642] <= 32'b11110100111101000000010111111000;
REG[6643] <= 32'b00000011000000001111110011110000;
REG[6644] <= 32'b11110000111111100000010111111101;
REG[6645] <= 32'b11111111111111110000111111100110;
REG[6646] <= 32'b11101100111111010000001111111100;
REG[6647] <= 32'b00000010111110110000001011110111;
REG[6648] <= 32'b11111011111100001111101000001011;
REG[6649] <= 32'b00000001111110001111101011101110;
REG[6650] <= 32'b11110101000000000000010011111100;
REG[6651] <= 32'b11111100111100101110111111111110;
REG[6652] <= 32'b00001101111111011111111011110111;
REG[6653] <= 32'b11110101000000110000010111111101;
REG[6654] <= 32'b00000010000000010010010000000011;
REG[6655] <= 32'b11110000111110001111110011110001;
REG[6656] <= 32'b00000101111111101111101000000011;
REG[6657] <= 32'b11111001111100111111100000000000;
REG[6658] <= 32'b00000100111111100001000100000000;
REG[6659] <= 32'b11111111111110010000001011111010;
REG[6660] <= 32'b11111111111101111111011011111101;
REG[6661] <= 32'b00010001111110111111110011101110;
REG[6662] <= 32'b11111111111111110000010111111000;
REG[6663] <= 32'b00001110111110010000000011111100;
REG[6664] <= 32'b11101110111111010000111000000100;
REG[6665] <= 32'b11110101111101001111100011111011;
REG[6666] <= 32'b00010011000011101111111100000001;
REG[6667] <= 32'b00000111000001100000000011111101;
REG[6668] <= 32'b11110100000001010000100100000011;
REG[6669] <= 32'b00100100000010001110111100001110;
REG[6670] <= 32'b00000001111111000010011000100000;
REG[6671] <= 32'b11110011000010011111100111111101;
REG[6672] <= 32'b11110111000011000000010100000100;
REG[6673] <= 32'b00000000111111111110110100000001;
REG[6674] <= 32'b11110110111111101111011100000101;
REG[6675] <= 32'b11110101000001100000001000000011;
REG[6676] <= 32'b00001100000011001111000111110100;
REG[6677] <= 32'b00000000111110010000011111111111;
REG[6678] <= 32'b11101110111101101111111000001001;
REG[6679] <= 32'b00100010000100001110111111110011;
REG[6680] <= 32'b11111011000000110000011000000000;
REG[6681] <= 32'b11101000111110000000111000000000;
REG[6682] <= 32'b11110011111110111111000011111011;
REG[6683] <= 32'b00001011111100111111110011110111;
REG[6684] <= 32'b11111111000001110000011100000010;
REG[6685] <= 32'b00010101111111111111100111100000;
REG[6686] <= 32'b00000000111111001111010111110100;
REG[6687] <= 32'b11110011111011010000011100000011;
REG[6688] <= 32'b11110100111101011111010111110001;
REG[6689] <= 32'b11110001000000011111101011111101;
REG[6690] <= 32'b00000110000001100000000100001001;
REG[6691] <= 32'b00010110000010011111110111111111;
REG[6692] <= 32'b11110100000101100001000011111000;
REG[6693] <= 32'b11111010000001010000010000010000;
REG[6694] <= 32'b11111111111101110000100111111001;
REG[6695] <= 32'b11110111111111010000001000000001;
REG[6696] <= 32'b00001110000000101111111011111101;
REG[6697] <= 32'b00000011000000000000001011111010;
REG[6698] <= 32'b11111011111110111111111100000000;
REG[6699] <= 32'b11111000111111000000000111111110;
REG[6700] <= 32'b00001000000101001111011011111000;
REG[6701] <= 32'b11111100111111000000011100000111;
REG[6702] <= 32'b11110110111110110000000111111011;
REG[6703] <= 32'b00000001000001001111010111111010;
REG[6704] <= 32'b00001100000010111110110111110001;
REG[6705] <= 32'b00000000111111000000100000001111;
REG[6706] <= 32'b11111000111101001111101111111100;
REG[6707] <= 32'b00000000000001101110111111101110;
REG[6708] <= 32'b11111101000010010000011011110010;
REG[6709] <= 32'b11101101111101111111000100000110;
REG[6710] <= 32'b00000010111110111111111000000110;
REG[6711] <= 32'b11111101000000110000001100001111;
REG[6712] <= 32'b00000010000010100000000100010001;
REG[6713] <= 32'b11101110111110000001000111110011;
REG[6714] <= 32'b00000011000110101111100011111111;
REG[6715] <= 32'b00101110000001010000010000000010;
REG[6716] <= 32'b11110101111101110000000011110100;
REG[6717] <= 32'b00010001001000100000100011111001;
REG[6718] <= 32'b11110001111100101111100100000000;
REG[6719] <= 32'b00001110000010100000110011111111;
REG[6720] <= 32'b00001000000010110000000111111111;
REG[6721] <= 32'b00010010000001101111001111101101;
REG[6722] <= 32'b00000110111110101111101111111001;
REG[6723] <= 32'b11110100111110000000110000000001;
REG[6724] <= 32'b00000111111110100000000011111100;
REG[6725] <= 32'b11111110000000000001000000010000;
REG[6726] <= 32'b11101111000000011111100000001001;
REG[6727] <= 32'b11111011111111011111001100001000;
REG[6728] <= 32'b11111100000001011111111000000010;
REG[6729] <= 32'b11110100000001111111110011110011;
REG[6730] <= 32'b11110010111101100000010000001001;
REG[6731] <= 32'b11111011000010000000001000000110;
REG[6732] <= 32'b11111111111111101111010000000101;
REG[6733] <= 32'b00001011000010101111100111110110;
REG[6734] <= 32'b11111001000000010000000000000100;
REG[6735] <= 32'b11111000000001010000111111111000;
REG[6736] <= 32'b00000111000001101111100000000000;
REG[6737] <= 32'b00001001000000011111001111101001;
REG[6738] <= 32'b11110010000001000000101111111110;
REG[6739] <= 32'b11110001111110010000101111111010;
REG[6740] <= 32'b11110110000010100000011100000101;
REG[6741] <= 32'b00000011111101010000000100000011;
REG[6742] <= 32'b00000111000001010001001100000100;
REG[6743] <= 32'b00000111111111110000011000000000;
REG[6744] <= 32'b11111111000010100001010000000111;
REG[6745] <= 32'b00000001111101101111011000000100;
REG[6746] <= 32'b00000011000001001111100111111011;
REG[6747] <= 32'b11111100000010010000011000000110;
REG[6748] <= 32'b11111100000100000000100011101111;
REG[6749] <= 32'b00000001111110101111101000010110;
REG[6750] <= 32'b00001000111100111111100011111010;
REG[6751] <= 32'b11111101000011010000011011110001;
REG[6752] <= 32'b11111111111110111111010011111100;
REG[6753] <= 32'b00001010000011010000011111110010;
REG[6754] <= 32'b11101010000000000000101000001101;
REG[6755] <= 32'b00000110111110001111110100001100;
REG[6756] <= 32'b00001100000100100000001100000101;
REG[6757] <= 32'b00000111000011001111001100000011;
REG[6758] <= 32'b00000001000001010000111100000001;
REG[6759] <= 32'b11110010111101001111110100000000;
REG[6760] <= 32'b00000100111110111111101100000011;
REG[6761] <= 32'b00000100000000100000010111111010;
REG[6762] <= 32'b11111100111101001111010100000000;
REG[6763] <= 32'b11111111000001001111101111111010;
REG[6764] <= 32'b11111100111101111111011111111111;
REG[6765] <= 32'b11111101111111101111110011110101;
REG[6766] <= 32'b11111100000001011111100111110011;
REG[6767] <= 32'b11110110111011001111011111110110;
REG[6768] <= 32'b11111101111101001111100111111011;
REG[6769] <= 32'b00010010000100101111101011110110;
REG[6770] <= 32'b11111100000000110000111100001011;
REG[6771] <= 32'b00000011111111100000000111110001;
REG[6772] <= 32'b11101101111100000000010111111001;
REG[6773] <= 32'b11110001111111101111100011110111;
REG[6774] <= 32'b11111101111111001111111111111010;
REG[6775] <= 32'b11111000111101000000011100000010;
REG[6776] <= 32'b11111100000010100000010100000111;
REG[6777] <= 32'b00010101000101111111011011111111;
REG[6778] <= 32'b00001000000100010000100100010101;
REG[6779] <= 32'b11111001111101110000011000010101;
REG[6780] <= 32'b11111001111110001111110100100010;
REG[6781] <= 32'b00001111111111101111100111111111;
REG[6782] <= 32'b00000000000110111111110111110010;
REG[6783] <= 32'b00000010000000011111100100001110;
REG[6784] <= 32'b11111110111101010000110000001010;
REG[6785] <= 32'b11101001000011110000110100010100;
REG[6786] <= 32'b00100001000111101110100100000101;
REG[6787] <= 32'b00000001000010100000111000010010;
REG[6788] <= 32'b00001100000001000001010000001010;
REG[6789] <= 32'b11111011111110100000011100010101;
REG[6790] <= 32'b11110110111100001111100011101111;
REG[6791] <= 32'b11111110111111101111101011110010;
REG[6792] <= 32'b11101101111100000000001100000000;
REG[6793] <= 32'b11110101111111111111110011111100;
REG[6794] <= 32'b00100001000000001111001111111110;
REG[6795] <= 32'b00000010000001010001010000000001;
REG[6796] <= 32'b11111000111011001111101000010001;
REG[6797] <= 32'b00011010000001001111111111101101;
REG[6798] <= 32'b00001110000011011111111011110010;
REG[6799] <= 32'b11111010111101100000100000010111;
REG[6800] <= 32'b00001111111101001111001100000001;
REG[6801] <= 32'b00010100000000111111110000100101;
REG[6802] <= 32'b00101011001101001111011011111001;
REG[6803] <= 32'b00011000000011100000100100001111;
REG[6804] <= 32'b11111010111110110001000000001100;
REG[6805] <= 32'b00001010000001100000000000000101;
REG[6806] <= 32'b00001001000001100000100000000100;
REG[6807] <= 32'b11111010000010010001001100000010;
REG[6808] <= 32'b00000110111101111111100100010001;
REG[6809] <= 32'b00010000000000001111100111101101;
REG[6810] <= 32'b00000001000101000000110111110101;
REG[6811] <= 32'b11110100111110011111101011111000;
REG[6812] <= 32'b00000101000000111111101111111111;
REG[6813] <= 32'b00000010111110111111111000000100;
REG[6814] <= 32'b11111101000000010000010100000100;
REG[6815] <= 32'b11111011000000101111101100000001;
REG[6816] <= 32'b00000100000010100000000011101100;
REG[6817] <= 32'b00001110000100100000000011111010;
REG[6818] <= 32'b11111011111011010011110000000001;
REG[6819] <= 32'b00000011000000000000000111101101;
REG[6820] <= 32'b11111010111101000000000011111101;
REG[6821] <= 32'b11111010111101110000001111111100;
REG[6822] <= 32'b11110001000001000000010111101010;
REG[6823] <= 32'b11111000111101111111001111111111;
REG[6824] <= 32'b00001011111101011111110011111111;
REG[6825] <= 32'b00000101111110101111000000010010;
REG[6826] <= 32'b11111101000010110000101000000011;
REG[6827] <= 32'b11111011000011111111011000000000;
REG[6828] <= 32'b11110111111010001111011111110111;
REG[6829] <= 32'b11111011000010000000011011110110;
REG[6830] <= 32'b11111110000001111111100000000100;
REG[6831] <= 32'b00110000000111110000100100100000;
REG[6832] <= 32'b11110101000101000000110000000010;
REG[6833] <= 32'b00001000111110001111110000000111;
REG[6834] <= 32'b00000010111111110000000011111110;
REG[6835] <= 32'b11110111111110001111100011111010;
REG[6836] <= 32'b11111000111111001111011111110101;
REG[6837] <= 32'b11111001111101101111100011110110;
REG[6838] <= 32'b11110000111010001111101100000001;
REG[6839] <= 32'b00001000000011110000110111111101;
REG[6840] <= 32'b11111101111110011111110100011110;
REG[6841] <= 32'b00100000111110100000000111110011;
REG[6842] <= 32'b00000001000101110001001011111111;
REG[6843] <= 32'b11101111111011101111011111111101;
REG[6844] <= 32'b11111111000011101111010011111100;
REG[6845] <= 32'b11111010111111011111011111111010;
REG[6846] <= 32'b11101101111110110000011011111101;
REG[6847] <= 32'b11101110111101101111011111110010;
REG[6848] <= 32'b00001001111110100000001000000011;
REG[6849] <= 32'b11111111111110010000100011111101;
REG[6850] <= 32'b00000111111101101111011111111010;
REG[6851] <= 32'b00001010000001000000111100000100;
REG[6852] <= 32'b00000100000101010000100011111100;
REG[6853] <= 32'b00000111000001010000011000010110;
REG[6854] <= 32'b00001000111111110000001100000010;
REG[6855] <= 32'b00000110111110101111001100001010;
REG[6856] <= 32'b00010101000001000000001011110010;
REG[6857] <= 32'b00000110111110011111111000001101;
REG[6858] <= 32'b00000000111100010000011111110001;
REG[6859] <= 32'b11110110000010000000011111111011;
REG[6860] <= 32'b00001101000010110000111100010000;
REG[6861] <= 32'b11110101000010100000010011111010;
REG[6862] <= 32'b11111111000001101110111100000001;
REG[6863] <= 32'b00010010000100010000101100000000;
REG[6864] <= 32'b11111100111110000001011100000100;
REG[6865] <= 32'b00000001000000111111011111101111;
REG[6866] <= 32'b11110001111100011111001011111101;
REG[6867] <= 32'b00000011000001011111111011101111;
REG[6868] <= 32'b11101011111011001111110111111100;
REG[6869] <= 32'b00000010111100111111100011110011;
REG[6870] <= 32'b11110111111110111111011011111001;
REG[6871] <= 32'b11111110111110101111101111111110;
REG[6872] <= 32'b11111101111100011111010111110001;
REG[6873] <= 32'b11111000111100011111000000000101;
REG[6874] <= 32'b11110101111100011111101011111110;
REG[6875] <= 32'b00000000111111010000111100000011;
REG[6876] <= 32'b11110101111100011111101100000111;
REG[6877] <= 32'b00010101000000001111101111110111;
REG[6878] <= 32'b00000110000001000000010111111100;
REG[6879] <= 32'b00000011111111111111110011111101;
REG[6880] <= 32'b00000111000010010000101100010000;
REG[6881] <= 32'b00000001111011000000000100000001;
REG[6882] <= 32'b00000011000011010000001011110111;
REG[6883] <= 32'b11111011111110011111100011111010;
REG[6884] <= 32'b00000011000011010000001100001000;
REG[6885] <= 32'b11111010111111110001001100010001;
REG[6886] <= 32'b00001011000000111111111011111110;
REG[6887] <= 32'b00000100000000101111110011111001;
REG[6888] <= 32'b11110110111101010000010000000000;
REG[6889] <= 32'b11111100111110101111011111110101;
REG[6890] <= 32'b11101111111110010000010000000100;
REG[6891] <= 32'b00000000111110111111101100001000;
REG[6892] <= 32'b11111000000001101111110011111100;
REG[6893] <= 32'b11110110111111110000111011110100;
REG[6894] <= 32'b11111000000101111111011111111100;
REG[6895] <= 32'b00001000111101011111011000000000;
REG[6896] <= 32'b11101111111110110000100011111001;
REG[6897] <= 32'b00000011000000101111010111110011;
REG[6898] <= 32'b00010100111111110001010000001011;
REG[6899] <= 32'b11110001111110100000011100000111;
REG[6900] <= 32'b00001000000100001111100111110100;
REG[6901] <= 32'b11111101000001111111001111110110;
REG[6902] <= 32'b11111100000000011111000011101110;
REG[6903] <= 32'b11110010111101010000000000011001;
REG[6904] <= 32'b00000011111100011111000111111010;
REG[6905] <= 32'b00001000000000110000010011110101;
REG[6906] <= 32'b11110101111011110000010100000101;
REG[6907] <= 32'b00010010000111101111001111101100;
REG[6908] <= 32'b11111010111110000000010000011000;
REG[6909] <= 32'b11111101111111001111111111111001;
REG[6910] <= 32'b11111001000010000001011100000101;
REG[6911] <= 32'b11111101111110001111011011111101;
REG[6912] <= 32'b00000111111110111111010100000000;
REG[6913] <= 32'b11111011111110111111110111111100;
REG[6914] <= 32'b00000010000010110000001011111100;
REG[6915] <= 32'b00010100000011000000000100000011;
REG[6916] <= 32'b00001011000100110001000100000101;
REG[6917] <= 32'b11111110111101001111110011111101;
REG[6918] <= 32'b00001001000001100000100011110111;
REG[6919] <= 32'b11111011000000111111110111111100;
REG[6920] <= 32'b11110100111100011111011111111110;
REG[6921] <= 32'b00000001111110001111000011111101;
REG[6922] <= 32'b11111101111110000000100011111101;
REG[6923] <= 32'b11110101111101001111001111110101;
REG[6924] <= 32'b00011011111111111111010111111010;
REG[6925] <= 32'b00000100111101010000011111110001;
REG[6926] <= 32'b11110111111110010000010011110011;
REG[6927] <= 32'b00001001000000100000001111111101;
REG[6928] <= 32'b00000101111110010000000011111101;
REG[6929] <= 32'b00000001000001010000101000000100;
REG[6930] <= 32'b11111110111111111111111000000110;
REG[6931] <= 32'b00001100000010100000000111101101;
REG[6932] <= 32'b11101110000101011111011100000100;
REG[6933] <= 32'b00000001000100110000101000001100;
REG[6934] <= 32'b00000100111111111111111100001111;
REG[6935] <= 32'b00001111000000001111111011111010;
REG[6936] <= 32'b11111101000101010001000111110100;
REG[6937] <= 32'b11111101111110010001000011111111;
REG[6938] <= 32'b00000000111111101111110111111010;
REG[6939] <= 32'b11111011111101001111110111110011;
REG[6940] <= 32'b11111110111110110000101100000001;
REG[6941] <= 32'b11111011111101101111010111111001;
REG[6942] <= 32'b11110001111111100000000100001110;
REG[6943] <= 32'b00000011000001010000110100011000;
REG[6944] <= 32'b00011100000011010001111100001001;
REG[6945] <= 32'b00001000000100100000100011110110;
REG[6946] <= 32'b00000011000001100001000011111100;
REG[6947] <= 32'b11110110000100001111001111110110;
REG[6948] <= 32'b00001011111111111111101100001110;
REG[6949] <= 32'b11101101000000010000001111111000;
REG[6950] <= 32'b11110111000000001110110011101101;
REG[6951] <= 32'b00000000000001111111111111101001;
REG[6952] <= 32'b00010000000010101111111000000011;
REG[6953] <= 32'b11111100111100110000110000000111;
REG[6954] <= 32'b11111101000010000000001011110101;
REG[6955] <= 32'b11111100111101011111111000000011;
REG[6956] <= 32'b00000110000101100001000100001001;
REG[6957] <= 32'b00000000000001110000010100010011;
REG[6958] <= 32'b00001110111110100000001000000110;
REG[6959] <= 32'b00000110000110000000001011110100;
REG[6960] <= 32'b11111000111101101111111011101100;
REG[6961] <= 32'b00000010111111011111011111111100;
REG[6962] <= 32'b11111111111110110000110100000011;
REG[6963] <= 32'b11110101000000000000000100001001;
REG[6964] <= 32'b00010110000010101111111011101001;
REG[6965] <= 32'b11110111111101101111110111110100;
REG[6966] <= 32'b00010000111101000000010011110100;
REG[6967] <= 32'b11111000111101001111010111101110;
REG[6968] <= 32'b11111101111111110000000111111100;
REG[6969] <= 32'b00001000111101101110101100000010;
REG[6970] <= 32'b11110010111111110001011000011011;
REG[6971] <= 32'b00011111001010101111110111111011;
REG[6972] <= 32'b00000101111101101111010100011110;
REG[6973] <= 32'b11111001111100001111100111110011;
REG[6974] <= 32'b11111000111110100001111000010101;
REG[6975] <= 32'b11110111111111010000010111111110;
REG[6976] <= 32'b00000101000000100000011011111111;
REG[6977] <= 32'b11110111111111000000001000000010;
REG[6978] <= 32'b00001100000000101111101111111010;
REG[6979] <= 32'b00000101000001111111100000000010;
REG[6980] <= 32'b00000100000001100000001100000101;
REG[6981] <= 32'b11111001111111000000001100010000;
REG[6982] <= 32'b00000010000000111111100011110111;
REG[6983] <= 32'b11110100000000111111101100001100;
REG[6984] <= 32'b00000111000000010000010011110111;
REG[6985] <= 32'b11110001111111000000001011111110;
REG[6986] <= 32'b11111111111110101111001000000010;
REG[6987] <= 32'b11110110111101101111010011101111;
REG[6988] <= 32'b11111001000001000000011100000100;
REG[6989] <= 32'b11110110111101000000010000001010;
REG[6990] <= 32'b00000101000001001111100011110011;
REG[6991] <= 32'b11111101000000010000101111111101;
REG[6992] <= 32'b11111110111111101111110011110100;
REG[6993] <= 32'b00000111000000110000000011110100;
REG[6994] <= 32'b11110100111110000000010011110110;
REG[6995] <= 32'b11110110000010011111110011110111;
REG[6996] <= 32'b00000110001000001111000011111011;
REG[6997] <= 32'b11111101111011100001010001001011;
REG[6998] <= 32'b11101000000100010001011011111101;
REG[6999] <= 32'b11110001111110111111010011111000;
REG[7000] <= 32'b11111010111011100000011011110011;
REG[7001] <= 32'b11111110000011110000111111110101;
REG[7002] <= 32'b11110101111110000000000011111111;
REG[7003] <= 32'b11111001111100111111110111110101;
REG[7004] <= 32'b11110111111110111111101111110101;
REG[7005] <= 32'b00001101000001000000001100000100;
REG[7006] <= 32'b11110111111110001111011011110101;
REG[7007] <= 32'b00010100000000110000010011111010;
REG[7008] <= 32'b00000000000000100001011100001110;
REG[7009] <= 32'b00011010000000101111100011110110;
REG[7010] <= 32'b11101001000010000000101100010010;
REG[7011] <= 32'b11111110000001111111101100001000;
REG[7012] <= 32'b11111101000011000000010100000100;
REG[7013] <= 32'b11110001000000011111110100000101;
REG[7014] <= 32'b11111011111101111111001111111100;
REG[7015] <= 32'b00000000111111011111100111101100;
REG[7016] <= 32'b11110010111110101111100011111111;
REG[7017] <= 32'b11111111111100011111101111111001;
REG[7018] <= 32'b11110111000000101110111011111101;
REG[7019] <= 32'b11111010111101001110100111110100;
REG[7020] <= 32'b11111100000000001111011011111010;
REG[7021] <= 32'b11111101000000101110001111101111;
REG[7022] <= 32'b11100110111111011111100000000100;
REG[7023] <= 32'b00000010000001110000001000000101;
REG[7024] <= 32'b00000101111111011111110100010000;
REG[7025] <= 32'b00010010000010000000101000000000;
REG[7026] <= 32'b00001000000010000001000111111110;
REG[7027] <= 32'b11111111111110111111110100000000;
REG[7028] <= 32'b11111100000001110000011000000011;
REG[7029] <= 32'b00000000000001000000000111111010;
REG[7030] <= 32'b11110100000001111111110100000000;
REG[7031] <= 32'b11110101000000011111011000000100;
REG[7032] <= 32'b11110110000000111111111111110011;
REG[7033] <= 32'b11111010000010111111101111110001;
REG[7034] <= 32'b11110101111011001111111100100100;
REG[7035] <= 32'b00001010111100100000001111101001;
REG[7036] <= 32'b00000000001000101111010011111111;
REG[7037] <= 32'b00000011000001100000000011111111;
REG[7038] <= 32'b11101010111011110001001000000010;
REG[7039] <= 32'b00000100111111001110111111101111;
REG[7040] <= 32'b00001101000011000000101100000000;
REG[7041] <= 32'b11111011111101111111010011111001;
REG[7042] <= 32'b00000011000000010001101000000101;
REG[7043] <= 32'b11110101000011010000101100000000;
REG[7044] <= 32'b00000111000001101111001000010001;
REG[7045] <= 32'b00000100111110101111101111110011;
REG[7046] <= 32'b11110011000000101111110100000101;
REG[7047] <= 32'b00000010111111001111111011111100;
REG[7048] <= 32'b11111001111111011111010011110010;
REG[7049] <= 32'b11110100000000101111101011111111;
REG[7050] <= 32'b11111101111110111111100000000011;
REG[7051] <= 32'b00000010111100010000011111111100;
REG[7052] <= 32'b11111111000010010000011100000001;
REG[7053] <= 32'b11111001000001101111010000001100;
REG[7054] <= 32'b00000011111111000000110100001000;
REG[7055] <= 32'b11100111000011001111100011111100;
REG[7056] <= 32'b00011011000110101111001100010100;
REG[7057] <= 32'b11111100111100000000000011111011;
REG[7058] <= 32'b11100100000010000000010111111000;
REG[7059] <= 32'b11111101111111011111101100000101;
REG[7060] <= 32'b11111000000000001111011000000110;
REG[7061] <= 32'b00000000111101101111011100000000;
REG[7062] <= 32'b11111100111110010000000100001100;
REG[7063] <= 32'b00000001111110110000110000001100;
REG[7064] <= 32'b00000100000000001111110100000011;
REG[7065] <= 32'b11111101000000010000000100000011;
REG[7066] <= 32'b11111001111111110001000000010110;
REG[7067] <= 32'b00011000000001111111011100000001;
REG[7068] <= 32'b00000001000000110000000100000001;
REG[7069] <= 32'b11111110111111001111110011111111;
REG[7070] <= 32'b00000111000001111111110011111010;
REG[7071] <= 32'b11111001111101100000101100001011;
REG[7072] <= 32'b00000000111110111111111111111100;
REG[7073] <= 32'b11111110000011110000011000001100;
REG[7074] <= 32'b11111001111110001111111000000011;
REG[7075] <= 32'b00010000000001001111101111110111;
REG[7076] <= 32'b11101100000010100000010011111111;
REG[7077] <= 32'b11111000000101101111110111111101;
REG[7078] <= 32'b11111001000010001111111000000110;
REG[7079] <= 32'b00001100111110011110111111111000;
REG[7080] <= 32'b11101110000100000000111011110000;
REG[7081] <= 32'b11110010111110100000000000000101;
REG[7082] <= 32'b11111100111111111111101100001011;
REG[7083] <= 32'b11110101111101111110101100000001;
REG[7084] <= 32'b00000000000001011111001111111110;
REG[7085] <= 32'b11101111000010110000111000001010;
REG[7086] <= 32'b00001010111110101111111100001101;
REG[7087] <= 32'b00011111000010001111111011111101;
REG[7088] <= 32'b00000011000010010000001100001011;
REG[7089] <= 32'b11110011111111001111101000001110;
REG[7090] <= 32'b11110101111110100000100011111001;
REG[7091] <= 32'b11110010000010110000011100001111;
REG[7092] <= 32'b00000011111110011110100100000000;
REG[7093] <= 32'b11111011000001000000000011111010;
REG[7094] <= 32'b11110001111111011111101000000000;
REG[7095] <= 32'b00000001111111011111000100000110;
REG[7096] <= 32'b11111100000000000000001011111111;
REG[7097] <= 32'b11110110000000110000000000000110;
REG[7098] <= 32'b00000100000000001111000000000111;
REG[7099] <= 32'b00000001000010001111101011110011;
REG[7100] <= 32'b11111100111110111111101000000000;
REG[7101] <= 32'b00001010111100001111100011110011;
REG[7102] <= 32'b11110101111101100000100111110001;
REG[7103] <= 32'b11110011111111001111100011111011;
REG[7104] <= 32'b00001111111111110000100100000101;
REG[7105] <= 32'b00000010111110100001000000000111;
REG[7106] <= 32'b00000110111111111111100111110001;
REG[7107] <= 32'b00000111111110110000010111110101;
REG[7108] <= 32'b11111101111110010000100100000111;
REG[7109] <= 32'b00000110111100011111001011110100;
REG[7110] <= 32'b11111001000001000000010111110010;
REG[7111] <= 32'b11110001111101011111000000001001;
REG[7112] <= 32'b00000011000000011111100111111011;
REG[7113] <= 32'b11110111111101110000001000001001;
REG[7114] <= 32'b11110111111101100000010011110110;
REG[7115] <= 32'b11111110111010011101010011001100;
REG[7116] <= 32'b11110001111100111111101000010011;
REG[7117] <= 32'b00000100111101101111100111110010;
REG[7118] <= 32'b11111100111111100000110100011110;
REG[7119] <= 32'b00010011000000011111010111110111;
REG[7120] <= 32'b11101101000010000000110011111001;
REG[7121] <= 32'b11110000000001011111100111111001;
REG[7122] <= 32'b11101110111010001111110100001100;
REG[7123] <= 32'b00011110000000010000110011110001;
REG[7124] <= 32'b00000000111111000000000111110100;
REG[7125] <= 32'b00011111111110101111100111111001;
REG[7126] <= 32'b11110100111100100000001100000100;
REG[7127] <= 32'b00001100111111011111011111111011;
REG[7128] <= 32'b00000111000010010001010111110110;
REG[7129] <= 32'b11110100111110000000011100010100;
REG[7130] <= 32'b00011101111101101111011011111001;
REG[7131] <= 32'b11100111111100011111001011110101;
REG[7132] <= 32'b11111011111101001111010011101101;
REG[7133] <= 32'b11101100111110111111001111110101;
REG[7134] <= 32'b11111100111110001111000100000010;
REG[7135] <= 32'b11110101111101110000100100000100;
REG[7136] <= 32'b11111011111101111111000011101111;
REG[7137] <= 32'b11111101111101101111010111110110;
REG[7138] <= 32'b11110111111110011111110100000010;
REG[7139] <= 32'b00000100111101011111110111111101;
REG[7140] <= 32'b11110000111010100001000100000011;
REG[7141] <= 32'b11101100111100001110110011100011;
REG[7142] <= 32'b00000111111010101111011011101110;
REG[7143] <= 32'b11111010111101100000111111110100;
REG[7144] <= 32'b00010011000000000001010000001100;
REG[7145] <= 32'b00001001000011011111100011110101;
REG[7146] <= 32'b11111000111110000000001000000011;
REG[7147] <= 32'b11110111111110000000011100000001;
REG[7148] <= 32'b00000111000000110000011011111010;
REG[7149] <= 32'b11111001111011111111110111110101;
REG[7150] <= 32'b11110111000001010000001011111001;
REG[7151] <= 32'b11111100111111101111011111111011;
REG[7152] <= 32'b00001010111101111111110100001010;
REG[7153] <= 32'b00011010111110110000101100001110;
REG[7154] <= 32'b00000010000010110001010000011000;
REG[7155] <= 32'b00000100000000010000101111101011;
REG[7156] <= 32'b11110000000001100000010100000000;
REG[7157] <= 32'b00000110111110100000010000001111;
REG[7158] <= 32'b11101101000000111111100100011011;
REG[7159] <= 32'b00010001000011001111010000001111;
REG[7160] <= 32'b11111101111110001111011111111000;
REG[7161] <= 32'b11110101111101111111011100000000;
REG[7162] <= 32'b00001000000000001111110011111010;
REG[7163] <= 32'b11110010111111001110100011101100;
REG[7164] <= 32'b11111111000010100000010111111111;
REG[7165] <= 32'b11111110000000001111110100000011;
REG[7166] <= 32'b00000001000000100000000000000100;
REG[7167] <= 32'b11110111111101111111111100000110;
REG[7168] <= 32'b00010100000001111111010011110110;
REG[7169] <= 32'b00000000111111001111111011111010;
REG[7170] <= 32'b11110101000000000000000100001101;
REG[7171] <= 32'b00000010000001011111010111111101;
REG[7172] <= 32'b11111110000001000000001011111100;
REG[7173] <= 32'b11110001111100111111100011111110;
REG[7174] <= 32'b11111110111111010000000011111100;
REG[7175] <= 32'b11110011111111101111101000001001;
REG[7176] <= 32'b11111000111111101111100100000001;
REG[7177] <= 32'b00010111111101101111110111110111;
REG[7178] <= 32'b00000110111101100000000011111100;
REG[7179] <= 32'b00010101000010100000101111110110;
REG[7180] <= 32'b00000011000000111111101100000100;
REG[7181] <= 32'b00011000000001101111010011111101;
REG[7182] <= 32'b11110101000001100001010111111011;
REG[7183] <= 32'b11101110111111111111100100001101;
REG[7184] <= 32'b00010110000011110000011011111111;
REG[7185] <= 32'b11111011111110001111111000010001;
REG[7186] <= 32'b00010001000011010000110111111111;
REG[7187] <= 32'b00000010111110010000011000001011;
REG[7188] <= 32'b00000001111110110000001100000001;
REG[7189] <= 32'b00000000111101110000100011111100;
REG[7190] <= 32'b00000101111101101111010111111110;
REG[7191] <= 32'b00000111111101101111111000000000;
REG[7192] <= 32'b00001110111111100000101000000000;
REG[7193] <= 32'b11111110000011100000010011110101;
REG[7194] <= 32'b00001000111011101101100011111110;
REG[7195] <= 32'b11111011111110100000100111110001;
REG[7196] <= 32'b11101110111110001110100111111001;
REG[7197] <= 32'b00000111111101101111001111111111;
REG[7198] <= 32'b11111101111111100000001011111110;
REG[7199] <= 32'b11111111111101011111111011111110;
REG[7200] <= 32'b00000110000000100000100111111010;
REG[7201] <= 32'b00001010000000110000010000001001;
REG[7202] <= 32'b00001110111111001111110011101010;
REG[7203] <= 32'b11100111000000010001001000000110;
REG[7204] <= 32'b00000110111111111111000111110110;
REG[7205] <= 32'b00010101111111101111101000000000;
REG[7206] <= 32'b11111010111111010001100011110111;
REG[7207] <= 32'b11110000111110011111101011111010;
REG[7208] <= 32'b00000001000000110000111000000111;
REG[7209] <= 32'b11111111000000100000010000000100;
REG[7210] <= 32'b00000100111111111111110111111100;
REG[7211] <= 32'b00000001000100010000110011111110;
REG[7212] <= 32'b00000101000000101111110000001010;
REG[7213] <= 32'b00000110000010101111111011110111;
REG[7214] <= 32'b11110110000001011111100000001011;
REG[7215] <= 32'b11111110111111101111110000000001;
REG[7216] <= 32'b11101001000010110000100011111011;
REG[7217] <= 32'b11110011000001101111111000000010;
REG[7218] <= 32'b00000011111110001111011100000101;
REG[7219] <= 32'b00000011111111000000010111111101;
REG[7220] <= 32'b11110000111111110000111000010111;
REG[7221] <= 32'b11110001111100100000100100010010;
REG[7222] <= 32'b00010000111111101110110011011101;
REG[7223] <= 32'b00000010111110100000001000001110;
REG[7224] <= 32'b11101111110111100000000100000011;
REG[7225] <= 32'b11111011000001001111101111110010;
REG[7226] <= 32'b11110101111101110000011000001011;
REG[7227] <= 32'b00001000000011010000001111111100;
REG[7228] <= 32'b00000100111110110000111100010100;
REG[7229] <= 32'b00000001111110110000010111111011;
REG[7230] <= 32'b00011000000010101111011100001000;
REG[7231] <= 32'b00000100000000110000001011111000;
REG[7232] <= 32'b11111101000000110000011011110000;
REG[7233] <= 32'b11111000111100011111001100010111;
REG[7234] <= 32'b00001011111110001111111111111000;
REG[7235] <= 32'b11111000111110001111010011110111;
REG[7236] <= 32'b00011011000010011111101111111010;
REG[7237] <= 32'b11110101111100110000100000000010;
REG[7238] <= 32'b11111000111111011111001111101110;
REG[7239] <= 32'b00001011111100000000001000010000;
REG[7240] <= 32'b00011101000010010001010011101111;
REG[7241] <= 32'b00000011000000111111111100000000;
REG[7242] <= 32'b00001100111101110000001000001000;
REG[7243] <= 32'b00001000111110000000010011110111;
REG[7244] <= 32'b11110011000000011111101011110011;
REG[7245] <= 32'b00001000000000111111101111110111;
REG[7246] <= 32'b11110000111101010000011000000011;
REG[7247] <= 32'b11111101111101011111001111111001;
REG[7248] <= 32'b11111101000001000000010111110110;
REG[7249] <= 32'b11110101111110001111111011111101;
REG[7250] <= 32'b00000001111111011111110111111111;
REG[7251] <= 32'b11110111111100011110110111111111;
REG[7252] <= 32'b00000100000001010000001000000000;
REG[7253] <= 32'b11111011111111111111110000000101;
REG[7254] <= 32'b11111111111101111111010011111100;
REG[7255] <= 32'b00000101000001101111110111110110;
REG[7256] <= 32'b11110111000100100001001000001100;
REG[7257] <= 32'b11111101000001001111101100000100;
REG[7258] <= 32'b00000001000011001110100011101110;
REG[7259] <= 32'b11110110111111001111111100000011;
REG[7260] <= 32'b11110000000000100001100100001001;
REG[7261] <= 32'b00001001000011011111110000001001;
REG[7262] <= 32'b11111110000000000000000100000000;
REG[7263] <= 32'b11110111000011010000100111110101;
REG[7264] <= 32'b11100001111000001111110111111001;
REG[7265] <= 32'b11101111000100001110011011110000;
REG[7266] <= 32'b11101101000000001111101111111001;
REG[7267] <= 32'b11110110000001011110100111110100;
REG[7268] <= 32'b11110101111110001111100000000011;
REG[7269] <= 32'b11101111111010011110111111111011;
REG[7270] <= 32'b11101110111111011111110100000001;
REG[7271] <= 32'b11111111000010110000011011110111;
REG[7272] <= 32'b11111100111111001111001111111001;
REG[7273] <= 32'b11110010111010011111111111111110;
REG[7274] <= 32'b11110100000000000001000011110110;
REG[7275] <= 32'b11110100111110001111010011110101;
REG[7276] <= 32'b11111000000001001111011100000010;
REG[7277] <= 32'b11111110111100001111010100000100;
REG[7278] <= 32'b11101001111101001110110011111100;
REG[7279] <= 32'b11110111000001000000000000000100;
REG[7280] <= 32'b00000000111111010000001011111110;
REG[7281] <= 32'b00000001000000101111101011111010;
REG[7282] <= 32'b11111000111110001111110000000110;
REG[7283] <= 32'b11110111000010000000001100000101;
REG[7284] <= 32'b11101110111011101111010100000010;
REG[7285] <= 32'b11111011000000110000000011101011;
REG[7286] <= 32'b11101110111111111111110000000001;
REG[7287] <= 32'b00011100000011010000000111111000;
REG[7288] <= 32'b11111010111111000001000000001011;
REG[7289] <= 32'b11101101111110100000000100010100;
REG[7290] <= 32'b00010001000111111110010111111010;
REG[7291] <= 32'b11101010000001011111001011111000;
REG[7292] <= 32'b11110010000000101110001000000001;
REG[7293] <= 32'b11111011111111011111111000000101;
REG[7294] <= 32'b00000010000010111110011011111011;
REG[7295] <= 32'b11111111111110111111101100000000;
REG[7296] <= 32'b00010011111110101111010100000011;
REG[7297] <= 32'b00000100000001110000010111111101;
REG[7298] <= 32'b11110110111111011111110000000001;
REG[7299] <= 32'b00011101000001111111011011111001;
REG[7300] <= 32'b00000000000001000000100100001111;
REG[7301] <= 32'b00000010111110110000111011110100;
REG[7302] <= 32'b00000000000011000000110111110010;
REG[7303] <= 32'b11111001111110101111010011111011;
REG[7304] <= 32'b00000011111100100000010100000000;
REG[7305] <= 32'b11111011111100111111001111111010;
REG[7306] <= 32'b00000000000000011111011000000010;
REG[7307] <= 32'b00010001111110011111100011110001;
REG[7308] <= 32'b00000110000011000000111100000000;
REG[7309] <= 32'b00010011000011001111101111111011;
REG[7310] <= 32'b00011010000000010001100100010101;
REG[7311] <= 32'b00001111000010110001000100010010;
REG[7312] <= 32'b00011000001000101111001111101101;
REG[7313] <= 32'b00000101000010010000110100010001;
REG[7314] <= 32'b11011110110111001111001011111101;
REG[7315] <= 32'b00000100000101010000101100000000;
REG[7316] <= 32'b11111011000011010000001011111001;
REG[7317] <= 32'b00001011000001101111011111110001;
REG[7318] <= 32'b11110110111010100000101000000100;
REG[7319] <= 32'b11110111111110011111101111110111;
REG[7320] <= 32'b11111111000100110000111100001111;
REG[7321] <= 32'b11111111000001011111011100000001;
REG[7322] <= 32'b00001011000000011111010111111001;
REG[7323] <= 32'b00011111000010010000001000001000;
REG[7324] <= 32'b11111001000000000000001011110010;
REG[7325] <= 32'b11111101111111110001001011111111;
REG[7326] <= 32'b00010100111110101111111111110011;
REG[7327] <= 32'b00001010000011100000011011111101;
REG[7328] <= 32'b00001000111101100001100000100000;
REG[7329] <= 32'b11110101111111111111111111111010;
REG[7330] <= 32'b00000101000001001111001011111100;
REG[7331] <= 32'b11111100111110101111101000000001;
REG[7332] <= 32'b00010111111101111111110000000001;
REG[7333] <= 32'b11111110000000100000101000000000;
REG[7334] <= 32'b11111011111110111111100000000001;
REG[7335] <= 32'b11111100111110001111010000000011;
REG[7336] <= 32'b11111001000011001111010011110101;
REG[7337] <= 32'b11110110000010000000011100000011;
REG[7338] <= 32'b00000001111111101111011111110100;
REG[7339] <= 32'b11110100111101011111101011110110;
REG[7340] <= 32'b11111001111101001111011111111001;
REG[7341] <= 32'b00100000000010001111010011111011;
REG[7342] <= 32'b11111010111110101111011111110001;
REG[7343] <= 32'b11110110111110000000111000000001;
REG[7344] <= 32'b00001011111111111111011011110111;
REG[7345] <= 32'b00000110000000100010001100010010;
REG[7346] <= 32'b11110101111010111111100111111111;
REG[7347] <= 32'b00000001000101000010001100000111;
REG[7348] <= 32'b11111111111111111111000111110110;
REG[7349] <= 32'b00011000000001111111111011111100;
REG[7350] <= 32'b11100100111000101110111100001100;
REG[7351] <= 32'b11110101111110001110110111110011;
REG[7352] <= 32'b11111110000011100000001000000000;
REG[7353] <= 32'b11101100111100111111110011111101;
REG[7354] <= 32'b00000011111111111111001011111110;
REG[7355] <= 32'b00000011000001010000000011110100;
REG[7356] <= 32'b00000110000001000000100000000000;
REG[7357] <= 32'b00001110000010001110111100000000;
REG[7358] <= 32'b00001001111101100000010100000101;
REG[7359] <= 32'b11100010111010010000001111101001;
REG[7360] <= 32'b00000000000010000001000111110111;
REG[7361] <= 32'b11110110000100001111100000000110;
REG[7362] <= 32'b00011100111101101111100100001000;
REG[7363] <= 32'b11111001111111010000100011110011;
REG[7364] <= 32'b11110001111011111111000011110110;
REG[7365] <= 32'b00011100000010000000001011110101;
REG[7366] <= 32'b00000011111110101111000111101011;
REG[7367] <= 32'b11101100111111010000010111110010;
REG[7368] <= 32'b11110010111100011111100111110010;
REG[7369] <= 32'b00000000111011011111000100000000;
REG[7370] <= 32'b00000011111100001111101100000110;
REG[7371] <= 32'b11110100000000101111101100000000;
REG[7372] <= 32'b11110101000000001111110000000011;
REG[7373] <= 32'b11101101111111111111101011110100;
REG[7374] <= 32'b00001001000000011111101111110000;
REG[7375] <= 32'b11111100000000101111110011110110;
REG[7376] <= 32'b11101000111110011111110011111110;
REG[7377] <= 32'b11101101111110001110111011111111;
REG[7378] <= 32'b00000111000000010000001011111100;
REG[7379] <= 32'b11110011111110010000000111110100;
REG[7380] <= 32'b11110011111101111110101000010000;
REG[7381] <= 32'b00010100111000001111010111110110;
REG[7382] <= 32'b11110100001001100001011111100111;
REG[7383] <= 32'b00010011000110010001010011111111;
REG[7384] <= 32'b11111000111110101111111111111110;
REG[7385] <= 32'b11110110111111000000000111111010;
REG[7386] <= 32'b11101110111011001110100111110010;
REG[7387] <= 32'b11111000111101110000001111111000;
REG[7388] <= 32'b11111010000000110000100011110100;
REG[7389] <= 32'b00000010111110011111010011111011;
REG[7390] <= 32'b11110001111011011111111111110110;
REG[7391] <= 32'b11111010111111001111110111111010;
REG[7392] <= 32'b00001101000100100000100011111001;
REG[7393] <= 32'b00000011111111110000110000000001;
REG[7394] <= 32'b11111001000000100000011111111001;
REG[7395] <= 32'b11111100111110011111000100000010;
REG[7396] <= 32'b00001011111101111111011111110111;
REG[7397] <= 32'b11110110111111111111010111110011;
REG[7398] <= 32'b11110100000001110000000000000011;
REG[7399] <= 32'b11111110111111101111010100001000;
REG[7400] <= 32'b00000011111111001111010111111000;
REG[7401] <= 32'b11110111111010001110101100001110;
REG[7402] <= 32'b00010110000011011111101011110010;
REG[7403] <= 32'b11101111000000001111111100001011;
REG[7404] <= 32'b00010110001000010001101000000100;
REG[7405] <= 32'b11110001000101010001110100001010;
REG[7406] <= 32'b00011101111110101111011111111110;
REG[7407] <= 32'b00001111000001100000000111111110;
REG[7408] <= 32'b00000101000001101110110011110100;
REG[7409] <= 32'b11111101111101111111110111111111;
REG[7410] <= 32'b11111011000010001111110100011001;
REG[7411] <= 32'b00001111000011001111111100000101;
REG[7412] <= 32'b00001100000100000000100100000000;
REG[7413] <= 32'b00000110000000100000011000000001;
REG[7414] <= 32'b00000010111110000000010100010010;
REG[7415] <= 32'b00011001111101011111010011111100;
REG[7416] <= 32'b11111011111111010000011011110110;
REG[7417] <= 32'b11110010111101001111100111110101;
REG[7418] <= 32'b00000101111110110001000000000111;
REG[7419] <= 32'b11111011111110011111011100000101;
REG[7420] <= 32'b11110110111110010000001100000101;
REG[7421] <= 32'b00000110111111111111010011111011;
REG[7422] <= 32'b11111011111111110000111111111001;
REG[7423] <= 32'b11111010111111010000001111111110;
REG[7424] <= 32'b11111101000011110001000100001000;
REG[7425] <= 32'b00000110000000110000001011111101;
REG[7426] <= 32'b00000000000000101111100011111000;
REG[7427] <= 32'b11111000000101110010001100010110;
REG[7428] <= 32'b11110111111011010000100000000110;
REG[7429] <= 32'b00000111111110011111010111111110;
REG[7430] <= 32'b11111110111101100001001111111111;
REG[7431] <= 32'b11111100000100111111010111110100;
REG[7432] <= 32'b00001000111100010000010100110100;
REG[7433] <= 32'b11011110111111001111010100001101;
REG[7434] <= 32'b11101110000101111110001111110111;
REG[7435] <= 32'b11110000000011001111001011110001;
REG[7436] <= 32'b11111000111110011111010100001100;
REG[7437] <= 32'b11110001000001101111110100000011;
REG[7438] <= 32'b00000101111100111111001000000101;
REG[7439] <= 32'b00001100111111001111111111111100;
REG[7440] <= 32'b00000001111111110000001100000110;
REG[7441] <= 32'b11111111000001000000011000010110;
REG[7442] <= 32'b00000011111101111111111111111011;
REG[7443] <= 32'b00000111000010010000111100000010;
REG[7444] <= 32'b00000010111101011111110000000101;
REG[7445] <= 32'b00000011000101010000100111110100;
REG[7446] <= 32'b11101111000100011111001111111110;
REG[7447] <= 32'b11110000111110000000001100000010;
REG[7448] <= 32'b11111111111100001111011011111111;
REG[7449] <= 32'b00001001000000110000011111110101;
REG[7450] <= 32'b11111010111110111111101011101100;
REG[7451] <= 32'b11101110111101111111001111110101;
REG[7452] <= 32'b00001110111110001111111100010011;
REG[7453] <= 32'b00001111000011100000001000000000;
REG[7454] <= 32'b00001001111110111110101111110111;
REG[7455] <= 32'b11101110111110100000100111111110;
REG[7456] <= 32'b11111101000001101110110111110111;
REG[7457] <= 32'b00000101000000111111101000000101;
REG[7458] <= 32'b00000111000100000000111100000001;
REG[7459] <= 32'b11111011000000100000000100010101;
REG[7460] <= 32'b00010000000111110001111100011001;
REG[7461] <= 32'b00010010000010000000101100000011;
REG[7462] <= 32'b00000111111110110000000100000110;
REG[7463] <= 32'b00000100000011010000100111111100;
REG[7464] <= 32'b11111001111110000000001000001010;
REG[7465] <= 32'b00010010111100110000001000001011;
REG[7466] <= 32'b00001100000100100000101100001001;
REG[7467] <= 32'b00000110000011100000100111111111;
REG[7468] <= 32'b00000001000010110000111100011010;
REG[7469] <= 32'b00000101111101101111010111110111;
REG[7470] <= 32'b00000110000101110001010111111110;
REG[7471] <= 32'b11110110111010101111111100001111;
REG[7472] <= 32'b00001101000100110001001111111101;
REG[7473] <= 32'b11111001111101010000010011110101;
REG[7474] <= 32'b11111110000010100000011000000101;
REG[7475] <= 32'b00001000111110001111100000000110;
REG[7476] <= 32'b00000110000001100000000000001110;
REG[7477] <= 32'b00000000000010000000001111110011;
REG[7478] <= 32'b00000000111101011110111111101010;
REG[7479] <= 32'b11111111111100101111011011110101;
REG[7480] <= 32'b11110100111011001111111111111011;
REG[7481] <= 32'b11111011111110011111011011110100;
REG[7482] <= 32'b00011100000011000000011011111100;
REG[7483] <= 32'b11111110111111100000011011111000;
REG[7484] <= 32'b00000001111111111111001011110111;
REG[7485] <= 32'b11111111111101111111110111111100;
REG[7486] <= 32'b11110011111110100000010111111011;
REG[7487] <= 32'b11111111111110101111100011101101;
REG[7488] <= 32'b11110110111101101111010111111000;
REG[7489] <= 32'b11111000111101011111010111111101;
REG[7490] <= 32'b11111011111110011111110111110001;
REG[7491] <= 32'b00000101111110100000001000000101;
REG[7492] <= 32'b00000111111110000001001011111100;
REG[7493] <= 32'b00001100000010100000000111111011;
REG[7494] <= 32'b00000010111111011111110000010010;
REG[7495] <= 32'b00001011000000000000110000000010;
REG[7496] <= 32'b11111110000011100000111000010111;
REG[7497] <= 32'b00001000111111001111011000000001;
REG[7498] <= 32'b11110010111101110000000100000001;
REG[7499] <= 32'b00000010000101110001010000011001;
REG[7500] <= 32'b11110110000000000000100100001101;
REG[7501] <= 32'b00010000000110001111111000001000;
REG[7502] <= 32'b11110100000011101111111000010100;
REG[7503] <= 32'b11111011111100111111010000001101;
REG[7504] <= 32'b11110001111111001111110000010011;
REG[7505] <= 32'b00010101000110100000101100001000;
REG[7506] <= 32'b00010111000100100000110100001111;
REG[7507] <= 32'b00000011111110110000010111111000;
REG[7508] <= 32'b00000111000100110000101100001011;
REG[7509] <= 32'b11111000000000101111101111111100;
REG[7510] <= 32'b11111110111111101110111011111100;
REG[7511] <= 32'b00000010000001011111110011111100;
REG[7512] <= 32'b11110010000001100000000000010000;
REG[7513] <= 32'b00001100000000000001100100000010;
REG[7514] <= 32'b11111010111100011111010011110101;
REG[7515] <= 32'b00000010000000011111110100010001;
REG[7516] <= 32'b00010110000000000000010100000111;
REG[7517] <= 32'b00001001000000011111111011110010;
REG[7518] <= 32'b11111100111101111110111111111110;
REG[7519] <= 32'b00000010000110010000000111111000;
REG[7520] <= 32'b11110100111111101111110100000101;
REG[7521] <= 32'b00001100000000100000011111110011;
REG[7522] <= 32'b11100111000101001110111111111010;
REG[7523] <= 32'b00011001111111011111110111110111;
REG[7524] <= 32'b11110100111111011111100111111011;
REG[7525] <= 32'b00000010111101010000001000001001;
REG[7526] <= 32'b11111011111101011111110011111001;
REG[7527] <= 32'b11110111000000010000010111111100;
REG[7528] <= 32'b00001001000010001111011011111111;
REG[7529] <= 32'b00000011000000000000100000000011;
REG[7530] <= 32'b11111111111111010000001111111011;
REG[7531] <= 32'b00000000111111001111111100000110;
REG[7532] <= 32'b11110110111110110000010111111000;
REG[7533] <= 32'b00000000111101101110110111111111;
REG[7534] <= 32'b00001110000001011111111111110100;
REG[7535] <= 32'b00000000111110111111011011111000;
REG[7536] <= 32'b00000111000001111111110111111001;
REG[7537] <= 32'b00000111000000110000000011111100;
REG[7538] <= 32'b11110111111101100001000011111101;
REG[7539] <= 32'b00000011111110111111010011110100;
REG[7540] <= 32'b00000010111101010000000011111001;
REG[7541] <= 32'b11111110111111101111100011110011;
REG[7542] <= 32'b11111111111111011111111100000010;
REG[7543] <= 32'b11111010111111010000000011110110;
REG[7544] <= 32'b11110100111111001111010011111011;
REG[7545] <= 32'b11101111000001010000101100000010;
REG[7546] <= 32'b11110101111101011110011111110101;
REG[7547] <= 32'b11111100111111111111101111111100;
REG[7548] <= 32'b11110101000000001111111111110101;
REG[7549] <= 32'b00000000000001000000001100010010;
REG[7550] <= 32'b00000010111111101111110100000010;
REG[7551] <= 32'b11111010000011010000010011111010;
REG[7552] <= 32'b11111010000001111111110100000000;
REG[7553] <= 32'b00000101111111100000100000001110;
REG[7554] <= 32'b11110100001001000001010000001000;
REG[7555] <= 32'b00000001111111111111001100101100;
REG[7556] <= 32'b01000010000010000000010100000110;
REG[7557] <= 32'b00000011000000110001101011111111;
REG[7558] <= 32'b11111011111111010000101011111111;
REG[7559] <= 32'b00000011111111110000011100000001;
REG[7560] <= 32'b00001101000011110000000011111111;
REG[7561] <= 32'b11111011000000000000100011111101;
REG[7562] <= 32'b11111001111110101111011111111011;
REG[7563] <= 32'b00000100111111101111010111111011;
REG[7564] <= 32'b00010111000011010000101000000110;
REG[7565] <= 32'b00000110111101110000101100000111;
REG[7566] <= 32'b00000110111111110000011100000010;
REG[7567] <= 32'b00001001000001100000001000001011;
REG[7568] <= 32'b11111011111110011111000111110011;
REG[7569] <= 32'b11111000000010111111110111111001;
REG[7570] <= 32'b11110101111011010000001100011001;
REG[7571] <= 32'b00001010111011011111000111101111;
REG[7572] <= 32'b11110100111111000000010011111001;
REG[7573] <= 32'b11111111000001011111010111110100;
REG[7574] <= 32'b11111011111110001111101100000001;
REG[7575] <= 32'b11110101111100111111100100001011;
REG[7576] <= 32'b00000110000011001111011000010100;
REG[7577] <= 32'b00000110111011001111010011101111;
REG[7578] <= 32'b11111001000111100001000111111011;
REG[7579] <= 32'b11111111111101000000000000001000;
REG[7580] <= 32'b00000100000011110000010111111110;
REG[7581] <= 32'b11111101111110100000011000000010;
REG[7582] <= 32'b00000000111111101111111011111101;
REG[7583] <= 32'b00001111000001100000011011111101;
REG[7584] <= 32'b00000000000000010000100100000111;
REG[7585] <= 32'b00000110111111111111101100001011;
REG[7586] <= 32'b00000000111110111111001111111111;
REG[7587] <= 32'b11110111000001010000011011111110;
REG[7588] <= 32'b11111111111111110000010011110101;
REG[7589] <= 32'b11111011000001110000101000001100;
REG[7590] <= 32'b00000111111111100000100011111111;
REG[7591] <= 32'b00000001111011110000011100001110;
REG[7592] <= 32'b00011001111110111111110111110111;
REG[7593] <= 32'b00001110000011000000100111111110;
REG[7594] <= 32'b11111100111111100001101000100010;
REG[7595] <= 32'b00010000111110010001000000000001;
REG[7596] <= 32'b00100100001100100010000100000100;
REG[7597] <= 32'b00000001111111000000111000001000;
REG[7598] <= 32'b11110011111110100000011011111101;
REG[7599] <= 32'b11110011000010001111011111110110;
REG[7600] <= 32'b11111101111110101111111100001100;
REG[7601] <= 32'b11111101000000010000111100000000;
REG[7602] <= 32'b11111101111111001111011011111000;
REG[7603] <= 32'b11111011111111010001010000000110;
REG[7604] <= 32'b00000000111101111111011111111001;
REG[7605] <= 32'b00000100111001001111000111110001;
REG[7606] <= 32'b11101001111011100001011011111100;
REG[7607] <= 32'b00000001111100101110100111111011;
REG[7608] <= 32'b11111111000000000000001111110011;
REG[7609] <= 32'b11110111111111000000011000010000;
REG[7610] <= 32'b11110101111010001111100100000010;
REG[7611] <= 32'b00000100000001011111001111101000;
REG[7612] <= 32'b11110001111111010000000011111101;
REG[7613] <= 32'b00001000000011001111110111110111;
REG[7614] <= 32'b00001110000100110000100100001000;
REG[7615] <= 32'b00001011111111100000001100000011;
REG[7616] <= 32'b11111000000001011111111111111001;
REG[7617] <= 32'b00010010000001010000001000000111;
REG[7618] <= 32'b00000001111111000000001111110011;
REG[7619] <= 32'b11111001000001001111101111111100;
REG[7620] <= 32'b00000010111110111111010000000001;
REG[7621] <= 32'b11111010111110000000010100001111;
REG[7622] <= 32'b00010010000000000000001000001011;
REG[7623] <= 32'b00000010000001100000001100000011;
REG[7624] <= 32'b00000000000001111111111100000010;
REG[7625] <= 32'b11111011000010001111111000000110;
REG[7626] <= 32'b11111010111111000000001100010100;
REG[7627] <= 32'b00001000111111011111110100000000;
REG[7628] <= 32'b00001000000100000000000111111101;
REG[7629] <= 32'b00000001000000100000010000001110;
REG[7630] <= 32'b00001010000000110000100111111101;
REG[7631] <= 32'b00010000000000000000011011111011;
REG[7632] <= 32'b00000111000000100001011011110011;
REG[7633] <= 32'b00000100111111011111110100000010;
REG[7634] <= 32'b00001110000000000000000000000011;
REG[7635] <= 32'b00001000111110011111001011111101;
REG[7636] <= 32'b00000111000011010000011011111001;
REG[7637] <= 32'b11111001111000101111010111111110;
REG[7638] <= 32'b11111111111111011111110111101000;
REG[7639] <= 32'b11111000000010001111110111111010;
REG[7640] <= 32'b11110101000010101111011111110001;
REG[7641] <= 32'b11111011111110001110111100001001;
REG[7642] <= 32'b00000000111100111111100100001011;
REG[7643] <= 32'b11111101000010010000010111111110;
REG[7644] <= 32'b11110011000001111111111011110110;
REG[7645] <= 32'b11110101111100011111000011111111;
REG[7646] <= 32'b11111000111110001111000111101110;
REG[7647] <= 32'b11101110111101000000010111111001;
REG[7648] <= 32'b11110101111100010000010000000110;
REG[7649] <= 32'b11110110111111010000001011101101;
REG[7650] <= 32'b00000011000100110000111000010001;
REG[7651] <= 32'b00111100000001010001001000001011;
REG[7652] <= 32'b00000111111111000001010011111000;
REG[7653] <= 32'b11111100111110111111001111111101;
REG[7654] <= 32'b11111001111110100000101000010010;
REG[7655] <= 32'b11110111111110111111011111111011;
REG[7656] <= 32'b00000110000100101111010011111110;
REG[7657] <= 32'b11110101111110100000110100001110;
REG[7658] <= 32'b00001101000000010000100111111100;
REG[7659] <= 32'b11111011000101000000101000001000;
REG[7660] <= 32'b00001011111111101111110100010111;
REG[7661] <= 32'b00000111000000110001011000000000;
REG[7662] <= 32'b11011111111100001111100000000001;
REG[7663] <= 32'b00000000111100011111001011110010;
REG[7664] <= 32'b11110101000010101111101011101111;
REG[7665] <= 32'b00000100000001111111001100000010;
REG[7666] <= 32'b11111000111011100000011011110101;
REG[7667] <= 32'b00001010111111111111010000000011;
REG[7668] <= 32'b00000000111111110000010011111010;
REG[7669] <= 32'b11101111000000000000001011111000;
REG[7670] <= 32'b00001011111111011111111100001101;
REG[7671] <= 32'b11111000000001010001000011101001;
REG[7672] <= 32'b11111011000010111111011000000011;
REG[7673] <= 32'b00010001111011101111001000000010;
REG[7674] <= 32'b00000000111111000000011011101111;
REG[7675] <= 32'b11110110000010100001010011111101;
REG[7676] <= 32'b00001001111100001111110111111000;
REG[7677] <= 32'b00010001111011100000100000000100;
REG[7678] <= 32'b00001100000000010001000111110111;
REG[7679] <= 32'b00000010000001100000000111111010;
REG[7680] <= 32'b11111000111110001110011011110100;
REG[7681] <= 32'b11101111111010111111100111110111;
REG[7682] <= 32'b11101100111110100000011111110100;
REG[7683] <= 32'b11110110111011001111000011111001;
REG[7684] <= 32'b11111011111011000000011000000111;
REG[7685] <= 32'b00000011111110111111011011110100;
REG[7686] <= 32'b00010110000100110000000011110110;
REG[7687] <= 32'b11111000111101100000111000010001;
REG[7688] <= 32'b11111011000001010000100100000001;
REG[7689] <= 32'b11111111111110110000001100000110;
REG[7690] <= 32'b00001011111111010000100011110110;
REG[7691] <= 32'b00000000000010000000101000001001;
REG[7692] <= 32'b11111000000000000000011100000010;
REG[7693] <= 32'b00001100000000110001100111111100;
REG[7694] <= 32'b11110100000011011111110111111011;
REG[7695] <= 32'b00001111111101101110110000011101;
REG[7696] <= 32'b11111010111101011111101100000000;
REG[7697] <= 32'b11111001001000100000001100000010;
REG[7698] <= 32'b11111000000000101111100111110101;
REG[7699] <= 32'b11111100111110111110110000000100;
REG[7700] <= 32'b11111110111110010000000111111111;
REG[7701] <= 32'b11110100000000110000000011110110;
REG[7702] <= 32'b11110110000000011111110100000001;
REG[7703] <= 32'b00001000000000001111011011111011;
REG[7704] <= 32'b11111010000000100000101111110011;
REG[7705] <= 32'b00000001000001111111110011111111;
REG[7706] <= 32'b00000001111100010000100000011000;
REG[7707] <= 32'b11111001111100011111101111110101;
REG[7708] <= 32'b11110100111101010000010011110111;
REG[7709] <= 32'b11111110000000011110110111110000;
REG[7710] <= 32'b11111100111111100000100011110100;
REG[7711] <= 32'b11110011111101111111111100000000;
REG[7712] <= 32'b00001001111101001111101100000000;
REG[7713] <= 32'b11111100111111110000000011110011;
REG[7714] <= 32'b11111000000010111111010011111000;
REG[7715] <= 32'b11111110111110001111011100000000;
REG[7716] <= 32'b00000110000101010000111111111101;
REG[7717] <= 32'b11111001111101011111110100000111;
REG[7718] <= 32'b00000011000011100000100011111111;
REG[7719] <= 32'b11111110111101000000000111111110;
REG[7720] <= 32'b11101010000000110000011011110000;
REG[7721] <= 32'b11111110111100011111101111111001;
REG[7722] <= 32'b11111110111100011111010100111001;
REG[7723] <= 32'b00011000111100101111110000001001;
REG[7724] <= 32'b00001101000110010000101011101110;
REG[7725] <= 32'b00000101000001001111100111111010;
REG[7726] <= 32'b00000001000001110000101100011000;
REG[7727] <= 32'b11110101000000100000000100000111;
REG[7728] <= 32'b00000111000011100000000111111111;
REG[7729] <= 32'b00001000000011011111101000000011;
REG[7730] <= 32'b00001100000100000000001011111111;
REG[7731] <= 32'b11110001111111110000100011111011;
REG[7732] <= 32'b11111100000000110001010100001100;
REG[7733] <= 32'b11111101000011100000101100000101;
REG[7734] <= 32'b11111010111101001111101111101110;
REG[7735] <= 32'b11100111111101110000011111110011;
REG[7736] <= 32'b11111101111100011110101111111010;
REG[7737] <= 32'b00000100111100111111001011110110;
REG[7738] <= 32'b11111011000000011111011011111000;
REG[7739] <= 32'b11111011111111011111110011111000;
REG[7740] <= 32'b11110110111111101111110011110011;
REG[7741] <= 32'b11111000111101111111000011110110;
REG[7742] <= 32'b00000100111110001111110011111001;
REG[7743] <= 32'b11111011000001110000110100001010;
REG[7744] <= 32'b00001000000001011111100011111100;
REG[7745] <= 32'b11111101000100010001000100001111;
REG[7746] <= 32'b00000001000000100000001000010101;
REG[7747] <= 32'b00000100000011101111100111110111;
REG[7748] <= 32'b11100111000101000000101000000001;
REG[7749] <= 32'b11101111111101001111001100001011;
REG[7750] <= 32'b00000011000000011111101111110000;
REG[7751] <= 32'b11101100000011011111111011110001;
REG[7752] <= 32'b11110011111111011111101111110000;
REG[7753] <= 32'b11110100000101111111001111110110;
REG[7754] <= 32'b11111100111111000000100011111011;
REG[7755] <= 32'b11111110111110101111101011110101;
REG[7756] <= 32'b11111100000100111111001011111100;
REG[7757] <= 32'b00001101000000101111001011110010;
REG[7758] <= 32'b11111001000001000001100100000001;
REG[7759] <= 32'b11110110000000100000001011111001;
REG[7760] <= 32'b00000111000000101111011111111100;
REG[7761] <= 32'b11110110111100111111110100100010;
REG[7762] <= 32'b00010111000010001111010111101110;
REG[7763] <= 32'b11110100111100101110001111111111;
REG[7764] <= 32'b11110010111011111111110111111000;
REG[7765] <= 32'b11110011000010010000001100000101;
REG[7766] <= 32'b00000101000101100000101000001010;
REG[7767] <= 32'b11111011000001111111111000010001;
REG[7768] <= 32'b00001010000011011111010111110111;
REG[7769] <= 32'b11111011111111011111101100000100;
REG[7770] <= 32'b00000001111110010000001011111001;
REG[7771] <= 32'b11111111000010111111001111110100;
REG[7772] <= 32'b11111010111100001111100100001001;
REG[7773] <= 32'b11111100111110011111110111111010;
REG[7774] <= 32'b00000111000100001111011100000001;
REG[7775] <= 32'b11111101111100101111101100000110;
REG[7776] <= 32'b11110111000000011111110111110100;
REG[7777] <= 32'b11110110111110010000001000000001;
REG[7778] <= 32'b11111111111111101111101111110110;
REG[7779] <= 32'b11110101111111111111111100000101;
REG[7780] <= 32'b11110011111111101111111000001000;
REG[7781] <= 32'b00000001000000001111010111111101;
REG[7782] <= 32'b11110111111111101111110011111010;
REG[7783] <= 32'b11110001111110000000000000001000;
REG[7784] <= 32'b00000100000011010000101100001100;
REG[7785] <= 32'b11111111000011000000100000001110;
REG[7786] <= 32'b11111111111111101111111100001101;
REG[7787] <= 32'b00010110000010001111001111111100;
REG[7788] <= 32'b00000100111111000000000000000100;
REG[7789] <= 32'b00000001000011111111101111101101;
REG[7790] <= 32'b11101110000110000001110000001101;
REG[7791] <= 32'b00000000000000100000011100011010;
REG[7792] <= 32'b00000110000011011111111000000100;
REG[7793] <= 32'b11110100000010011111111011110000;
REG[7794] <= 32'b11110110111111110000010100001010;
REG[7795] <= 32'b11111111111110000000000111111011;
REG[7796] <= 32'b11110110000010011111110111110101;
REG[7797] <= 32'b00000110111110111111100111111110;
REG[7798] <= 32'b11110101111100000000100111111101;
REG[7799] <= 32'b11110110000101001111110100000001;
REG[7800] <= 32'b00000010111100111111011100000011;
REG[7801] <= 32'b11110010000000110000011000000001;
REG[7802] <= 32'b00000000111110110000010000001101;
REG[7803] <= 32'b00000000000000000000010011101100;
REG[7804] <= 32'b11111001000000100000100100001111;
REG[7805] <= 32'b00001100111101101111111111111010;
REG[7806] <= 32'b11111100000000001111100011111111;
REG[7807] <= 32'b00001001000001110000100100001001;
REG[7808] <= 32'b11110011111011001111001011111011;
REG[7809] <= 32'b11110100111101011111111000000001;
REG[7810] <= 32'b00001011000000100001110000001010;
REG[7811] <= 32'b11111010000011000000010000010000;
REG[7812] <= 32'b00000010111111111111110100000001;
REG[7813] <= 32'b00000000000000100000000011110001;
REG[7814] <= 32'b11110010000000001111100111111000;
REG[7815] <= 32'b11110111111101111111001011110000;
REG[7816] <= 32'b11110100111101111111110000000001;
REG[7817] <= 32'b11110111111101001111011011111100;
REG[7818] <= 32'b11111110000000001111111100000110;
REG[7819] <= 32'b11110110000000011111110011111010;
REG[7820] <= 32'b00000011111110010000000111110101;
REG[7821] <= 32'b00000000000001011111110111110101;
REG[7822] <= 32'b11111101111111111111101011110110;
REG[7823] <= 32'b11110110111110000000000000001001;
REG[7824] <= 32'b11111011111110011111111111111010;
REG[7825] <= 32'b00010010111110110000011000000111;
REG[7826] <= 32'b11111101000001110010111100000110;
REG[7827] <= 32'b00000010000001110000101111110110;
REG[7828] <= 32'b11111100111101001111111111111010;
REG[7829] <= 32'b11110011111110110000011100010011;
REG[7830] <= 32'b00000010111110011111000011111100;
REG[7831] <= 32'b11111011000011111111110100000100;
REG[7832] <= 32'b00000000000000111111100000001000;
REG[7833] <= 32'b00001001001100100000011000000100;
REG[7834] <= 32'b11111010000000111111110000000000;
REG[7835] <= 32'b11110100000101001111101011111011;
REG[7836] <= 32'b00010000111110001111001111111011;
REG[7837] <= 32'b00000010000010100000001100001010;
REG[7838] <= 32'b00000110111011011111010011101100;
REG[7839] <= 32'b00010000000011001111111011111101;
REG[7840] <= 32'b11111001111100110000010111111110;
REG[7841] <= 32'b11111000111011111111010111110111;
REG[7842] <= 32'b11111011111100011110110111111110;
REG[7843] <= 32'b11110111111101011111111111111001;
REG[7844] <= 32'b11110100000001011111110111111100;
REG[7845] <= 32'b00001011111111001111010100000010;
REG[7846] <= 32'b11111101111101110000001011111110;
REG[7847] <= 32'b00000010111111101111110011111011;
REG[7848] <= 32'b00000101000010010000111111111110;
REG[7849] <= 32'b00000111000011010000001000001111;
REG[7850] <= 32'b00000110111101100000001000001111;
REG[7851] <= 32'b11111010111101001110110011111010;
REG[7852] <= 32'b00000110000010101111111011110100;
REG[7853] <= 32'b11101010111110110000100000000000;
REG[7854] <= 32'b00010110000010101110110111101110;
REG[7855] <= 32'b11110111000000010000000100010001;
REG[7856] <= 32'b00011110111111100000000100000011;
REG[7857] <= 32'b11111100000010000001100011111110;
REG[7858] <= 32'b00001110000100001111101011111111;
REG[7859] <= 32'b00000101111110000001010100010101;
REG[7860] <= 32'b00001000111111110001011011110100;
REG[7861] <= 32'b11110100000001001111110011110111;
REG[7862] <= 32'b00000100111011101110101100000010;
REG[7863] <= 32'b00000000000010010000111011111010;
REG[7864] <= 32'b11110110000011110000010011111110;
REG[7865] <= 32'b11101010111010110000001100000011;
REG[7866] <= 32'b00000110000010101111000111111001;
REG[7867] <= 32'b00001100000000011111100111111101;
REG[7868] <= 32'b00000101111111000000101000000101;
REG[7869] <= 32'b11111101111011110000111100000101;
REG[7870] <= 32'b00000010111110001111101111110000;
REG[7871] <= 32'b11111111111111100000011011111101;
REG[7872] <= 32'b00000001111100111111001111111000;
REG[7873] <= 32'b11111111111111110001010100001001;
REG[7874] <= 32'b11111111000010111111011011110111;
REG[7875] <= 32'b00000111000011000000010100010011;
REG[7876] <= 32'b00110010000010110000001000000010;
REG[7877] <= 32'b11111110111101000001010011111101;
REG[7878] <= 32'b11111010111110001111011011111100;
REG[7879] <= 32'b00000110111111001111110111111111;
REG[7880] <= 32'b11111101000000010001001000000000;
REG[7881] <= 32'b11101111111101000000000000000000;
REG[7882] <= 32'b00000101000000100001011000010011;
REG[7883] <= 32'b00000110111111011111011000000001;
REG[7884] <= 32'b00001111000110010001001000000011;
REG[7885] <= 32'b11111100000000011111010100000001;
REG[7886] <= 32'b00001100111111111111111000000001;
REG[7887] <= 32'b00000010000000111111001011111110;
REG[7888] <= 32'b00001001000001100000010011110111;
REG[7889] <= 32'b11110010111110100000000100000001;
REG[7890] <= 32'b00000011000000011111010000000011;
REG[7891] <= 32'b00000101000010101111111011111110;
REG[7892] <= 32'b00000010111111010000000011111011;
REG[7893] <= 32'b00000111000000110000001100000111;
REG[7894] <= 32'b00001111000011100000100100001011;
REG[7895] <= 32'b00000110111111010000011000000100;
REG[7896] <= 32'b00000001111101110000111011101011;
REG[7897] <= 32'b11101111111110000001010111111010;
REG[7898] <= 32'b11111011111100001111111100001100;
REG[7899] <= 32'b00011100000100111111101111111011;
REG[7900] <= 32'b11110011000011010000000000001001;
REG[7901] <= 32'b11111110000010010000111000001100;
REG[7902] <= 32'b00010110000011101111010000001110;
REG[7903] <= 32'b00001010000100110000100011111110;
REG[7904] <= 32'b11111001000001111111111111111110;
REG[7905] <= 32'b11111110000001100000101100001100;
REG[7906] <= 32'b00000011111110111111011000000011;
REG[7907] <= 32'b00010110000000101111010011111101;
REG[7908] <= 32'b00000011000011010010001100000100;
REG[7909] <= 32'b11111000000000110001110000010010;
REG[7910] <= 32'b11110000000001100000010100000110;
REG[7911] <= 32'b00100101000111011110000100000110;
REG[7912] <= 32'b00000101111111100001100000000110;
REG[7913] <= 32'b11101011000110100000001111110011;
REG[7914] <= 32'b00000011111111101111100000010000;
REG[7915] <= 32'b00010010111010100000110100001100;
REG[7916] <= 32'b11111010000101000000111111101010;
REG[7917] <= 32'b11111001111110001111011100001111;
REG[7918] <= 32'b00001001111011000000101100000000;
REG[7919] <= 32'b11111010000001100000010100010010;
REG[7920] <= 32'b00010010000011101111101100000100;
REG[7921] <= 32'b11111111111110110000000011111100;
REG[7922] <= 32'b11110010000001110000001111111000;
REG[7923] <= 32'b11110101111110100000001111111100;
REG[7924] <= 32'b11111100000000111111010011110110;
REG[7925] <= 32'b00000001111100011111100111111101;
REG[7926] <= 32'b11101110111010001111011111111001;
REG[7927] <= 32'b11111011111111100000011100001010;
REG[7928] <= 32'b11111010000001101111101100000001;
REG[7929] <= 32'b11111111000001111111111000001010;
REG[7930] <= 32'b11111010111110011111100011111000;
REG[7931] <= 32'b11111100000001010000000011111000;
REG[7932] <= 32'b00010000111110010000101100000010;
REG[7933] <= 32'b00000010111110000001110011111101;
REG[7934] <= 32'b00000001111110001111111011101100;
REG[7935] <= 32'b00010010000100111111101011110111;
REG[7936] <= 32'b11111000111100100001000100000000;
REG[7937] <= 32'b11111010000101011111110011111100;
REG[7938] <= 32'b00001000000001000000001100001100;
REG[7939] <= 32'b11111111111111101111100000001000;
REG[7940] <= 32'b00001010111110011111010011111001;
REG[7941] <= 32'b00001000001010000010000000000001;
REG[7942] <= 32'b11110111000001011111011111111000;
REG[7943] <= 32'b00001110111111111111111100000011;
REG[7944] <= 32'b00000011111101111111010000000010;
REG[7945] <= 32'b11111011000010111111010111111111;
REG[7946] <= 32'b00001000000000001111110011110111;
REG[7947] <= 32'b11111011111110010000110111111110;
REG[7948] <= 32'b11111011000000001111111111111111;
REG[7949] <= 32'b00001110111111001111110011111100;
REG[7950] <= 32'b00010101000101101111001000001100;
REG[7951] <= 32'b00001100111101100000011100010111;
REG[7952] <= 32'b11111111111110011111111111110001;
REG[7953] <= 32'b11111100000011101111000011111001;
REG[7954] <= 32'b11111100111110100000101100001010;
REG[7955] <= 32'b00000000000001010000011011101010;
REG[7956] <= 32'b00000110000100000000010000000111;
REG[7957] <= 32'b00010010111101010000010000001011;
REG[7958] <= 32'b11111000000100110001111000000010;
REG[7959] <= 32'b00001011000001001111100000001111;
REG[7960] <= 32'b00000100111110000001111000000111;
REG[7961] <= 32'b11110011000101010000011011111111;
REG[7962] <= 32'b00001010000010001111100000001111;
REG[7963] <= 32'b00000010111111010000000000000110;
REG[7964] <= 32'b11111000000010100000000100001100;
REG[7965] <= 32'b11110111111111111111101000001010;
REG[7966] <= 32'b00001110111111101111110111111110;
REG[7967] <= 32'b11110101000001010001100000001000;
REG[7968] <= 32'b11111001000010110000100111111110;
REG[7969] <= 32'b00000111111101101111010100001001;
REG[7970] <= 32'b00001011000001000001110100010000;
REG[7971] <= 32'b00000101000011000000001000000101;
REG[7972] <= 32'b00010100000010001111000100000000;
REG[7973] <= 32'b00100101111111100000010000001010;
REG[7974] <= 32'b11110110001000000010100011111001;
REG[7975] <= 32'b11111111000001111111001111110001;
REG[7976] <= 32'b11111011000001000000100100000110;
REG[7977] <= 32'b00000011111111001111111111111100;
REG[7978] <= 32'b00000001111111010011001000000000;
REG[7979] <= 32'b00000101111111010000111000000100;
REG[7980] <= 32'b11111100111101011111101011100010;
REG[7981] <= 32'b11110111111111010001100011110101;
REG[7982] <= 32'b11111011000011011111111000000010;
REG[7983] <= 32'b00010010111010101111100100011010;
REG[7984] <= 32'b00010010000111101111110011111100;
REG[7985] <= 32'b00000100000011011111010011111001;
REG[7986] <= 32'b11110011111110001111101100000001;
REG[7987] <= 32'b11111110000001011111111011111010;
REG[7988] <= 32'b00000111000000111111101000001000;
REG[7989] <= 32'b00000000111101110000000000001010;
REG[7990] <= 32'b00001001000100011110111011111001;
REG[7991] <= 32'b11110110000001010000100000010111;
REG[7992] <= 32'b11110111111111101111010100011100;
REG[7993] <= 32'b00101110000111101111111100000110;
REG[7994] <= 32'b11111100001000000001110100011101;
REG[7995] <= 32'b11101010111110010000001011111001;
REG[7996] <= 32'b11110110111110011111010111111011;
REG[7997] <= 32'b11111001111110101111111000000000;
REG[7998] <= 32'b11110001111110001111100111111111;
REG[7999] <= 32'b00000010111110111111110100000110;
REG[8000] <= 32'b00011011111101100000000000000010;
REG[8001] <= 32'b00000001111111000001001011110001;
REG[8002] <= 32'b11111111000000001111100100000000;
REG[8003] <= 32'b00000110111101111111110111111011;
REG[8004] <= 32'b11111110000001100000111011111001;
REG[8005] <= 32'b11111101111110101111101100000111;
REG[8006] <= 32'b00001010111101001111011011111111;
REG[8007] <= 32'b00000110111111100000011011110111;
REG[8008] <= 32'b11111011000001101111111101001001;
REG[8009] <= 32'b00001010111110010000010111111011;
REG[8010] <= 32'b11111001000111101111010100000001;
REG[8011] <= 32'b00000000000000010000010100001010;
REG[8012] <= 32'b11101111000001101111111111111111;
REG[8013] <= 32'b11110010111101100000110111111000;
REG[8014] <= 32'b11110101111101011111101011111010;
REG[8015] <= 32'b11111110111011111111111011111000;
REG[8016] <= 32'b11110111111110100000001111110101;
REG[8017] <= 32'b11111100111101110000100100001011;
REG[8018] <= 32'b00001011111111100000001111111111;
REG[8019] <= 32'b00000111111111000000100111111001;
REG[8020] <= 32'b00000111111110010001000100001110;
REG[8021] <= 32'b00000101111110001111111011110100;
REG[8022] <= 32'b00001111000011010000000100000001;
REG[8023] <= 32'b00000101111111000001100000001001;
REG[8024] <= 32'b11110011000000000000110000001000;
REG[8025] <= 32'b00000110000100101111101100000000;
REG[8026] <= 32'b00001011000101100000000100001011;
REG[8027] <= 32'b00001110111111110001010100010001;
REG[8028] <= 32'b00001100000000110000101000000110;
REG[8029] <= 32'b00001110000010011111011000000101;
REG[8030] <= 32'b11111011111110100001000000000010;
REG[8031] <= 32'b00011011000011010001011111111111;
REG[8032] <= 32'b11111110111101000000110100010011;
REG[8033] <= 32'b00010010000000100000010111111110;
REG[8034] <= 32'b00010000000101000000110000000111;
REG[8035] <= 32'b00000110111111010000100011111000;
REG[8036] <= 32'b00000110000000001111101011111100;
REG[8037] <= 32'b00001000111110100000011000001000;
REG[8038] <= 32'b11111100111100110000001011110110;
REG[8039] <= 32'b00001000000001011111101111111010;
REG[8040] <= 32'b11111000111110111111101111111101;
REG[8041] <= 32'b11111101111010110000100100010111;
REG[8042] <= 32'b11111001111100110000100011110100;
REG[8043] <= 32'b11110110111110001111011111110011;
REG[8044] <= 32'b11110100111010101111011000000011;
REG[8045] <= 32'b00000101111110100000010000011011;
REG[8046] <= 32'b11111000000000010000011100000000;
REG[8047] <= 32'b00000010000110111111100100000011;
REG[8048] <= 32'b11111110000000011111010100001111;
REG[8049] <= 32'b11110011111111010000110111101110;
REG[8050] <= 32'b11110011000001101111001111111000;
REG[8051] <= 32'b00001010111011001111001111111110;
REG[8052] <= 32'b00000011000010010001011111111010;
REG[8053] <= 32'b11110100111111100001100111111101;
REG[8054] <= 32'b11110111000000100000010100000011;
REG[8055] <= 32'b00001000111111111110100000000100;
REG[8056] <= 32'b00000111000001110000000100000000;
REG[8057] <= 32'b11101101000001101111111011111100;
REG[8058] <= 32'b11101101111101001111011111111011;
REG[8059] <= 32'b11111001111111001111000011110101;
REG[8060] <= 32'b11110110111101011111110011111001;
REG[8061] <= 32'b11110100111111011111101111101111;
REG[8062] <= 32'b11111010111111001111100011110111;
REG[8063] <= 32'b11111010111101111111100011111011;
REG[8064] <= 32'b00001110111111001111101111111111;
REG[8065] <= 32'b00001000000010010001001000001101;
REG[8066] <= 32'b11111010000000011111101100000010;
REG[8067] <= 32'b00001010000001011111101011111111;
REG[8068] <= 32'b11110110111101010000100100000111;
REG[8069] <= 32'b11111111111111001111100111111101;
REG[8070] <= 32'b11111110000001011111100100001010;
REG[8071] <= 32'b00001011000010000000100011110101;
REG[8072] <= 32'b11111010000010011111010011111001;
REG[8073] <= 32'b11111001000000001111101011111101;
REG[8074] <= 32'b11101111111100000000000100001000;
REG[8075] <= 32'b00001000000000011111100011110111;
REG[8076] <= 32'b11111110111111001111101100000000;
REG[8077] <= 32'b11111001111110100001000100010010;
REG[8078] <= 32'b11110101111111001111101011111001;
REG[8079] <= 32'b11111011111111001110111100000101;
REG[8080] <= 32'b11111101111110111111101100001001;
REG[8081] <= 32'b11111111000011101111011011111011;
REG[8082] <= 32'b11111111000011100000010000010000;
REG[8083] <= 32'b00000100111100110000010000000110;
REG[8084] <= 32'b00000111000101110000100011111011;
REG[8085] <= 32'b00000101111111100001001000001000;
REG[8086] <= 32'b00000000111111110000000111110110;
REG[8087] <= 32'b00011101111111101111001111111010;
REG[8088] <= 32'b00001001000000110010000000000101;
REG[8089] <= 32'b11111001111111110000001111110111;
REG[8090] <= 32'b00000100111110011111101111111110;
REG[8091] <= 32'b00000010111111110001001011111101;
REG[8092] <= 32'b11111100111101100000000011111111;
REG[8093] <= 32'b00001110111110101111101111110111;
REG[8094] <= 32'b00000010000101000001000111110101;
REG[8095] <= 32'b11110110000000000000000100011111;
REG[8096] <= 32'b00101011000000011111011111111111;
REG[8097] <= 32'b00000001000011100000111011111110;
REG[8098] <= 32'b11110110111110000000110011111000;
REG[8099] <= 32'b11110111000010110001110100000010;
REG[8100] <= 32'b00000010111110111111010011111010;
REG[8101] <= 32'b00001010111101000000011111111010;
REG[8102] <= 32'b00000100000001100001000111110010;
REG[8103] <= 32'b00001110000100010000000100000000;
REG[8104] <= 32'b11110111111110101111110100010000;
REG[8105] <= 32'b00000100000001101111111111111000;
REG[8106] <= 32'b00000011000000100000001100000101;
REG[8107] <= 32'b11111001111101110000011111111011;
REG[8108] <= 32'b11111001000000110000110100000001;
REG[8109] <= 32'b00000010111010111111001100000000;
REG[8110] <= 32'b00000111000000110000001011111001;
REG[8111] <= 32'b11111101000001110000100000001100;
REG[8112] <= 32'b11111101000000001111111011110110;
REG[8113] <= 32'b00000001111111011111000000000101;
REG[8114] <= 32'b11111111000100100000111100010100;
REG[8115] <= 32'b11101101000010010000001011111100;
REG[8116] <= 32'b11110000111110101111110111111100;
REG[8117] <= 32'b00000000111110111111011111110111;
REG[8118] <= 32'b11111011000011000000000111111100;
REG[8119] <= 32'b11111111111101111111000100001011;
REG[8120] <= 32'b11110001111111011111100111111001;
REG[8121] <= 32'b11101110111010101111001100011100;
REG[8122] <= 32'b00001101000011000000000011110001;
REG[8123] <= 32'b11110000000000100000000111111101;
REG[8124] <= 32'b00000010111100101111100011101011;
REG[8125] <= 32'b11111100000000111110111111100001;
REG[8126] <= 32'b11100111111100001110011011101110;
REG[8127] <= 32'b00010000000000101110101111101111;
REG[8128] <= 32'b11101001111011000000011011111101;
REG[8129] <= 32'b11111001111010101110011111110001;
REG[8130] <= 32'b11111000111111110000000000000101;
REG[8131] <= 32'b11111101111111111111000111110001;
REG[8132] <= 32'b11110100111101011111001011111101;
REG[8133] <= 32'b11110111111101101111011011111001;
REG[8134] <= 32'b11111100000001010000110100001101;
REG[8135] <= 32'b00001101111110001111001100000010;
REG[8136] <= 32'b00000000000001101111011011110000;
REG[8137] <= 32'b11110001111111001111101100001111;
REG[8138] <= 32'b11111111111010101110100111110011;
REG[8139] <= 32'b11101111111100101111010100000110;
REG[8140] <= 32'b11111011111101101110100011101001;
REG[8141] <= 32'b11110000111101111111100011111000;
REG[8142] <= 32'b11110000111101001111001100000001;
REG[8143] <= 32'b00000100000010001111111011110001;
REG[8144] <= 32'b11110110111110001111111100000101;
REG[8145] <= 32'b11111000111110011111110011111100;
REG[8146] <= 32'b11111100111111111111001011110000;
REG[8147] <= 32'b11110111111111100000000011111101;
REG[8148] <= 32'b00000010111111010000100000000011;
REG[8149] <= 32'b00000110000000101110101111101111;
REG[8150] <= 32'b00010010111110111111011000000010;
REG[8151] <= 32'b00001001111111000000101000000000;
REG[8152] <= 32'b11110001000000011111101011111000;
REG[8153] <= 32'b00000110000010110000100100000001;
REG[8154] <= 32'b11110101111101010001001011111101;
REG[8155] <= 32'b00000100000010001111101100000111;
REG[8156] <= 32'b00010110111111111111011011111110;
REG[8157] <= 32'b00000010111100011110110111111011;
REG[8158] <= 32'b11111101000010101111110100000101;
REG[8159] <= 32'b00001101111101001111000000001001;
REG[8160] <= 32'b11110000000000100001000111111011;
REG[8161] <= 32'b11101100111101101111110000000001;
REG[8162] <= 32'b00000110111100111111111011111110;
REG[8163] <= 32'b11110111111110101111110000000001;
REG[8164] <= 32'b00010001000000011111110011111000;
REG[8165] <= 32'b11111111111110110000011011111100;
REG[8166] <= 32'b00000101000100110001001111111111;
REG[8167] <= 32'b00000110000001100000011000011000;
REG[8168] <= 32'b00011001111101010000000100000010;
REG[8169] <= 32'b11110010000000100000010011111110;
REG[8170] <= 32'b11110100111101111111010000000000;
REG[8171] <= 32'b11111110000001000000111000011001;
REG[8172] <= 32'b11111110001101010011001000001111;
REG[8173] <= 32'b00010101000001101111111100010011;
REG[8174] <= 32'b00100100000011011111110011110000;
REG[8175] <= 32'b11101110111100011111010111111100;
REG[8176] <= 32'b11111001000000111111000011110000;
REG[8177] <= 32'b11110011111101011111011000000101;
REG[8178] <= 32'b00000000111100101111011011110100;
REG[8179] <= 32'b11110100111111100000000011111011;
REG[8180] <= 32'b11111011111010111110101011110011;
REG[8181] <= 32'b00000010111101000000000111110011;
REG[8182] <= 32'b11101011111101000000101000000101;
REG[8183] <= 32'b00000110111100111110110111110011;
REG[8184] <= 32'b11110101000001111111001000000111;
REG[8185] <= 32'b00000101000001011111000000000010;
REG[8186] <= 32'b11111000111110110000011000000000;
REG[8187] <= 32'b11110111000011011111011011111001;
REG[8188] <= 32'b00000001111110101111010111111101;
REG[8189] <= 32'b11111111000010000001001100001000;
REG[8190] <= 32'b11101101111111110000010100010100;
REG[8191] <= 32'b00001111000000001110011011111111;
REG[8192] <= 32'b00000010000000100000000100000010;
REG[8193] <= 32'b11110100111110110000001000000001;
REG[8194] <= 32'b11111111000010101111101111111110;
REG[8195] <= 32'b11111101000000001111011000000111;
REG[8196] <= 32'b00001011000001011111010011111100;
REG[8197] <= 32'b11110100000001010000101011111111;
REG[8198] <= 32'b11111011000000010000001000001010;
REG[8199] <= 32'b00001101000011101111010111110111;
REG[8200] <= 32'b11110011111111100000111100010111;
REG[8201] <= 32'b11110101000001100000010011111110;
REG[8202] <= 32'b00010011000101110000101111111100;
REG[8203] <= 32'b11100110111010101111110100001111;
REG[8204] <= 32'b00000010000011001111100111101101;
REG[8205] <= 32'b11110011000011100000011000001010;
REG[8206] <= 32'b11111001111110110000110011111011;
REG[8207] <= 32'b11111100111110000000010100000110;
REG[8208] <= 32'b11111011111100010000001000011001;
REG[8209] <= 32'b00100111000110111110110011101011;
REG[8210] <= 32'b11111111000000000000011000000000;
REG[8211] <= 32'b00000111000010001111010000000111;
REG[8212] <= 32'b11111110000010000000011000011000;
REG[8213] <= 32'b00000111111111111111101111111011;
REG[8214] <= 32'b11111111000010000000100000000010;
REG[8215] <= 32'b00001101000111111111110111111100;
REG[8216] <= 32'b11111000000001011111110111111100;
REG[8217] <= 32'b00000100111101011111011100000000;
REG[8218] <= 32'b11111011000010000000011011111000;
REG[8219] <= 32'b11101111000001011111111100000011;
REG[8220] <= 32'b11111001111110101111110011111011;
REG[8221] <= 32'b00000001000010111111011111110100;
REG[8222] <= 32'b00001011000000000001001111111111;
REG[8223] <= 32'b00000011000010000001010111110101;
REG[8224] <= 32'b11111110111111000000101111111111;
REG[8225] <= 32'b11110101111100000000000000010111;
REG[8226] <= 32'b00000000111110011111001111101100;
REG[8227] <= 32'b11111101000100011111111111101101;
REG[8228] <= 32'b11110100111111000000011100000101;
REG[8229] <= 32'b00000000001000011110111100011001;
REG[8230] <= 32'b00001100000000001110100101000110;
REG[8231] <= 32'b11110000000101100001001000001101;
REG[8232] <= 32'b11110101000111100001001100000101;
REG[8233] <= 32'b00000101111110010000000111111101;
REG[8234] <= 32'b00000000000010000000000111101111;
REG[8235] <= 32'b00000110111100001111101100001100;
REG[8236] <= 32'b00010100111101100000011011110110;
REG[8237] <= 32'b11111010111111110000001111111111;
REG[8238] <= 32'b11111100111110001111011011111000;
REG[8239] <= 32'b00000101000100111111011111111011;
REG[8240] <= 32'b11110100111101111111111000000011;
REG[8241] <= 32'b00000011111111111110100000000010;
REG[8242] <= 32'b11111101000001111111110111110010;
REG[8243] <= 32'b11100110000010010000010011111010;
REG[8244] <= 32'b00000101111110111111111011111100;
REG[8245] <= 32'b11111111111100110000010100001000;
REG[8246] <= 32'b00011111111110001111111111110111;
REG[8247] <= 32'b11111100111110111111011011111011;
REG[8248] <= 32'b11111000111110000000010011111000;
REG[8249] <= 32'b11111001111110101111011011101010;
REG[8250] <= 32'b11111110111101111111110111111110;
REG[8251] <= 32'b11111101111101100000001111111110;
REG[8252] <= 32'b11101010000000101111011111111100;
REG[8253] <= 32'b11111101000000111111110011111001;
REG[8254] <= 32'b11101111111110101111100100001000;
REG[8255] <= 32'b11111101111100111110111111111000;
REG[8256] <= 32'b00001010111101101111001111111010;
REG[8257] <= 32'b00001000111100011111011111101001;
REG[8258] <= 32'b11100110111111011111110011100111;
REG[8259] <= 32'b00000011111101011111000011111000;
REG[8260] <= 32'b11110110111110101111000111110111;
REG[8261] <= 32'b11111111111111000000001111111100;
REG[8262] <= 32'b11111110000011010000111000000110;
REG[8263] <= 32'b00001001000000100000011000010101;
REG[8264] <= 32'b00010000000010010001000100000101;
REG[8265] <= 32'b11110101000000101111101100000010;
REG[8266] <= 32'b11111110111111000000000011110110;
REG[8267] <= 32'b00000000111111001111110111111111;
REG[8268] <= 32'b11111100000010010000000111111011;
REG[8269] <= 32'b00000110000001101110100000001101;
REG[8270] <= 32'b00010010000101110000001000001110;
REG[8271] <= 32'b11100110111100001101111000000010;
REG[8272] <= 32'b11110111111111000011011000010110;
REG[8273] <= 32'b00000001111101111111011011110000;
REG[8274] <= 32'b00000100000001011111110011111101;
REG[8275] <= 32'b00001000000110111111111100001010;
REG[8276] <= 32'b11111011111100100000000100000011;
REG[8277] <= 32'b11111010000010011111100111110001;
REG[8278] <= 32'b11110110111011110010010000100011;
REG[8279] <= 32'b00101001111111000000101000001011;
REG[8280] <= 32'b00001010000010010000111000000100;
REG[8281] <= 32'b00001101111111010000000000000010;
REG[8282] <= 32'b00000011111010111111010111111110;
REG[8283] <= 32'b11111101111110010000001111110101;
REG[8284] <= 32'b00000000000100110000010111111110;
REG[8285] <= 32'b11110100111111110000010000001011;
REG[8286] <= 32'b11110101111011011110111011111100;
REG[8287] <= 32'b00000000111111101111111011110001;
REG[8288] <= 32'b11110101111010101111111111111011;
REG[8289] <= 32'b11101011111001111111100111111111;
REG[8290] <= 32'b00001100000001100000001011110000;
REG[8291] <= 32'b11110110111110010000011100000100;
REG[8292] <= 32'b11110111111011101111101100000110;
REG[8293] <= 32'b11101110110111000000011011110110;
REG[8294] <= 32'b11111111111111111111011111110011;
REG[8295] <= 32'b11110001111101110000111000001000;
REG[8296] <= 32'b00000101000001011111010111111101;
REG[8297] <= 32'b11101011111110111111000100001101;
REG[8298] <= 32'b11110000001001101111111011110110;
REG[8299] <= 32'b11110011000011011111110100010001;
REG[8300] <= 32'b00010010000000000000000000001110;
REG[8301] <= 32'b11111101111100001111110011111100;
REG[8302] <= 32'b11111000000000010000010100000000;
REG[8303] <= 32'b11101110000000110001011000000000;
REG[8304] <= 32'b11101011111101101111000111111000;
REG[8305] <= 32'b11110001111111100001000100000110;
REG[8306] <= 32'b00000100111011001111011011111011;
REG[8307] <= 32'b00001000111111000000000111111001;
REG[8308] <= 32'b00000011111110000000010111111111;
REG[8309] <= 32'b11111110000010010000011011111000;
REG[8310] <= 32'b00000010111111101111110111111100;
REG[8311] <= 32'b11111001111110000000000000000000;
REG[8312] <= 32'b00000000111011101110110011110000;
REG[8313] <= 32'b11111110111111100000010111110111;
REG[8314] <= 32'b11110111111111001111110011111100;
REG[8315] <= 32'b11110100111110110011011100010111;
REG[8316] <= 32'b00000100000000010000000111110010;
REG[8317] <= 32'b00011110000001110001000000000010;
REG[8318] <= 32'b00001000110111101111010011110110;
REG[8319] <= 32'b11110111111110110000001000011000;
REG[8320] <= 32'b00010111000101001111111000000000;
REG[8321] <= 32'b00000110000101010000111100001101;
REG[8322] <= 32'b11111000000000110000010000001111;
REG[8323] <= 32'b00000101000010011110111011110111;
REG[8324] <= 32'b11111101000000100000110011110000;
REG[8325] <= 32'b11101100111011001111001111111010;
REG[8326] <= 32'b00000001111101011110011111110100;
REG[8327] <= 32'b11110111111111001111101011110111;
REG[8328] <= 32'b11111110111100111111011000001000;
REG[8329] <= 32'b00000101111111111111111111101011;
REG[8330] <= 32'b11101001111110111111011111110111;
REG[8331] <= 32'b11110110111011001111010111111011;
REG[8332] <= 32'b11111011111111000001110100001110;
REG[8333] <= 32'b00001101000000110000101111110001;
REG[8334] <= 32'b11111101111111100000100100010111;
REG[8335] <= 32'b00011110000001111111001100000101;
REG[8336] <= 32'b00000100000010010000100100000100;
REG[8337] <= 32'b00010100000010001111101000100111;
REG[8338] <= 32'b00001111111100001111101011111010;
REG[8339] <= 32'b11101100111111110000000111110000;
REG[8340] <= 32'b11101101000000010000101111110011;
REG[8341] <= 32'b11111100111110100000111100001111;
REG[8342] <= 32'b00001011000011000001001000000000;
REG[8343] <= 32'b00001000000001110000011000001101;
REG[8344] <= 32'b00011001111100011111111100000011;
REG[8345] <= 32'b00000000000000000000010111111000;
REG[8346] <= 32'b11111101111110111110101011111011;
REG[8347] <= 32'b00000000111111111111110111110101;
REG[8348] <= 32'b11101110111111110000001000000001;
REG[8349] <= 32'b11111100111100001111001000010001;
REG[8350] <= 32'b00001101000000011111011100000101;
REG[8351] <= 32'b11110010111110011111011111101111;
REG[8352] <= 32'b11110110000110000000110111110111;
REG[8353] <= 32'b11111011111100100000000100000100;
REG[8354] <= 32'b00010101111100101111001011110011;
REG[8355] <= 32'b11110011111010111110101100000000;
REG[8356] <= 32'b00000000111110101110111111101100;
REG[8357] <= 32'b11101010111111110000010011111101;
REG[8358] <= 32'b11101000111010111110011100000010;
REG[8359] <= 32'b00000100111111101111111100000100;
REG[8360] <= 32'b00000111111101010000100100000011;
REG[8361] <= 32'b00000001111101101111101111110011;
REG[8362] <= 32'b11111111111111010000001111111111;
REG[8363] <= 32'b11110100111011001111101100000100;
REG[8364] <= 32'b11111010111101101111111111111101;
REG[8365] <= 32'b11111010111101111111001111110001;
REG[8366] <= 32'b11110111000101100000000111111101;
REG[8367] <= 32'b00000010111110000000010000011000;
REG[8368] <= 32'b00000010111111100000011100001001;
REG[8369] <= 32'b00010011111101011110011111111000;
REG[8370] <= 32'b00000110000001010000110011101100;
REG[8371] <= 32'b11110011111101110000100100001000;
REG[8372] <= 32'b11111100111100011111111111111101;
REG[8373] <= 32'b11111101111100111110111011111010;
REG[8374] <= 32'b11111100111111111111100011101110;
REG[8375] <= 32'b11101010000001001111011000000001;
REG[8376] <= 32'b11111001111011111111001000001001;
REG[8377] <= 32'b00001001000110000000100100000101;
REG[8378] <= 32'b11111101000010001111011011101011;
REG[8379] <= 32'b00000000111110101111001100001111;
REG[8380] <= 32'b11110011111100110001101100010010;
REG[8381] <= 32'b11101100000011001111011111101001;
REG[8382] <= 32'b00000111000010001111001000001110;
REG[8383] <= 32'b11110100111101010000111100010010;
REG[8384] <= 32'b11101110000001111111010011110011;
REG[8385] <= 32'b00000111000010011111010000001001;
REG[8386] <= 32'b00000001111110010000011011111111;
REG[8387] <= 32'b11111100000010010001001111111011;
REG[8388] <= 32'b00000000111110111111110011111110;
REG[8389] <= 32'b00001000111110011111011111111101;
REG[8390] <= 32'b00010100111111001111010111110011;
REG[8391] <= 32'b00010010000110101111001111110100;
REG[8392] <= 32'b00001111000011010000111100100110;
REG[8393] <= 32'b11110100000011010000000100001011;
REG[8394] <= 32'b00010000000010111110111000000111;
REG[8395] <= 32'b11101110111101101111110111110010;
REG[8396] <= 32'b11110110111101001111011111101101;
REG[8397] <= 32'b00001001111101111111101011111101;
REG[8398] <= 32'b11111100111011110000110000000111;
REG[8399] <= 32'b00000011111111101111110011110110;
REG[8400] <= 32'b11110111111010111111010000001011;
REG[8401] <= 32'b00000000000001101111001011110010;
REG[8402] <= 32'b11111100000001100000100000001000;
REG[8403] <= 32'b11101100111010000000111000000100;
REG[8404] <= 32'b00001010111111111111100011111000;
REG[8405] <= 32'b11111110111100111110110111110111;
REG[8406] <= 32'b11111010111100011111010111101011;
REG[8407] <= 32'b11101111111001010000101000000110;
REG[8408] <= 32'b00001100111111001110111011111000;
REG[8409] <= 32'b11101010111101111111101100000000;
REG[8410] <= 32'b11101110111100010001010011111100;
REG[8411] <= 32'b11101010000110001111100111110001;
REG[8412] <= 32'b00001001111110101111100111111000;
REG[8413] <= 32'b11110111111100111111000111110000;
REG[8414] <= 32'b11111011111111000000100000001101;
REG[8415] <= 32'b11110101111100011111001111111111;
REG[8416] <= 32'b00001111000110011111100111111100;
REG[8417] <= 32'b11111110000010001111111000000001;
REG[8418] <= 32'b11110100111101111110111000000001;
REG[8419] <= 32'b11111111111101110000110111111110;
REG[8420] <= 32'b11110110000010000000001011111111;
REG[8421] <= 32'b00001101111100111111111000000101;
REG[8422] <= 32'b11111111111110010000001000001100;
REG[8423] <= 32'b11111111000010001111111100001100;
REG[8424] <= 32'b11111100001100000000011000001011;
REG[8425] <= 32'b11111001000010011111110000010101;
REG[8426] <= 32'b00000000111111111111110000000010;
REG[8427] <= 32'b00000000111101111111100011111110;
REG[8428] <= 32'b00001011000011110000011111111010;
REG[8429] <= 32'b11111000000000010000101000000001;
REG[8430] <= 32'b00000111111110111111011100000110;
REG[8431] <= 32'b11111111111110101111010111111001;
REG[8432] <= 32'b11111111111111010001001100010111;
REG[8433] <= 32'b11111101111111011111110011111000;
REG[8434] <= 32'b00010011000010001111100111111011;
REG[8435] <= 32'b11111010111100100000001100000000;
REG[8436] <= 32'b11110110111111000000001011111010;
REG[8437] <= 32'b11110110000001101110011100001011;
REG[8438] <= 32'b00010101000000001111001000001000;
REG[8439] <= 32'b00000001111110000000010000010010;
REG[8440] <= 32'b00000001000101001110101111100011;
REG[8441] <= 32'b11110010000010000001010100000000;
REG[8442] <= 32'b11101011111001011111000100001100;
REG[8443] <= 32'b00001110111110011111111111111000;
REG[8444] <= 32'b00000010111011001111100011111101;
REG[8445] <= 32'b00000000111110111111110111111111;
REG[8446] <= 32'b11110101111101011110110111111010;
REG[8447] <= 32'b11111111000011110000101011110111;
REG[8448] <= 32'b11110010111111010000010000001110;
REG[8449] <= 32'b00010011111110011110110111111010;
REG[8450] <= 32'b11110110000001110000011111111111;
REG[8451] <= 32'b11111000000001001111011011111111;
REG[8452] <= 32'b00000101000010010000000000000001;
REG[8453] <= 32'b11111011000001000000010100001010;
REG[8454] <= 32'b00010010000010101111110111101010;
REG[8455] <= 32'b11110011111011010000100111110111;
REG[8456] <= 32'b11110101111011011111010011101110;
REG[8457] <= 32'b11111001111111011111011011110100;
REG[8458] <= 32'b11111000111011011110010011111101;
REG[8459] <= 32'b11111001111111111111101011111000;
REG[8460] <= 32'b11110110000000001111111111110101;
REG[8461] <= 32'b11110111111100111111001111110011;
REG[8462] <= 32'b11100110000000011111010111111011;
REG[8463] <= 32'b00000001111111001111101100000000;
REG[8464] <= 32'b11111111111111110000101111110110;
REG[8465] <= 32'b11111010111111111111110111111100;
REG[8466] <= 32'b00001010111101000000000000000000;
REG[8467] <= 32'b00000010000000100001101000001100;
REG[8468] <= 32'b00000011000001010000001000000010;
REG[8469] <= 32'b00001011000000111110110111111001;
REG[8470] <= 32'b11111010000001111111110111110110;
REG[8471] <= 32'b11101111000010010001000100000101;
REG[8472] <= 32'b11111110111110011111010111101000;
REG[8473] <= 32'b11110111111000000000010011111001;
REG[8474] <= 32'b00010011000000000011011111110011;
REG[8475] <= 32'b11111011111101100000110111101011;
REG[8476] <= 32'b11111001111011010000001000000011;
REG[8477] <= 32'b00000101111011001111101000000011;
REG[8478] <= 32'b11111100111110101111101111100111;
REG[8479] <= 32'b11101011111100001111011100000010;
REG[8480] <= 32'b00001101111100111111001011110110;
REG[8481] <= 32'b11111000000000100001010000001001;
REG[8482] <= 32'b11111010111110011111110100001101;
REG[8483] <= 32'b00001001000000111111001100000100;
REG[8484] <= 32'b00000100000110110001010100000011;
REG[8485] <= 32'b11111111111111101111110011111101;
REG[8486] <= 32'b11111110111111001111111111111110;
REG[8487] <= 32'b11111010111111000000000100010001;
REG[8488] <= 32'b00001110111101111111101011101100;
REG[8489] <= 32'b00000100000010110000011111111110;
REG[8490] <= 32'b00010100000000001110110000001110;
REG[8491] <= 32'b00001110000010010000011100011000;
REG[8492] <= 32'b11111111000011000001111000010001;
REG[8493] <= 32'b11111000111110100000011100000011;
REG[8494] <= 32'b00001011000010000000101100000111;
REG[8495] <= 32'b11111101111111100000010100000101;
REG[8496] <= 32'b00000101000011011111010111110000;
REG[8497] <= 32'b11101000111110111111110000000110;
REG[8498] <= 32'b11111100000001000000000000001000;
REG[8499] <= 32'b11110010111110000000001100000111;
REG[8500] <= 32'b00010101000011011111010111110111;
REG[8501] <= 32'b00001100111111100000011111111111;
REG[8502] <= 32'b11101010111100110001001111110101;
REG[8503] <= 32'b00000110111111100000110100010000;
REG[8504] <= 32'b00000110111111110000000000001000;
REG[8505] <= 32'b00000101000011100000011011101011;
REG[8506] <= 32'b11110000111101001111100011111111;
REG[8507] <= 32'b11110000111111000000001100000010;
REG[8508] <= 32'b00000101000011010000001111110101;
REG[8509] <= 32'b11101101111110110000010000010100;
REG[8510] <= 32'b00000001111111111110111111111000;
REG[8511] <= 32'b00000010000000100000011011110010;
REG[8512] <= 32'b11101111111110011111101111110100;
REG[8513] <= 32'b00000000111111110000011000000010;
REG[8514] <= 32'b11110101111100001111011000010100;
REG[8515] <= 32'b00011000000000001110101111101001;
REG[8516] <= 32'b11110010111111000001111000000110;
REG[8517] <= 32'b11111100000000011111101100000100;
REG[8518] <= 32'b00000100000001001111110011111110;
REG[8519] <= 32'b11110110000000001111111100001110;
REG[8520] <= 32'b00000001000000101111100100001010;
REG[8521] <= 32'b00001001000100101111111011110010;
REG[8522] <= 32'b11110101000011100001010100010011;
REG[8523] <= 32'b11111010111011101111100000000010;
REG[8524] <= 32'b00000000000001111111111111110100;
REG[8525] <= 32'b11101110111110100000000000001111;
REG[8526] <= 32'b00000010111100101110010100000010;
REG[8527] <= 32'b11111101000101011111100111110010;
REG[8528] <= 32'b11101111111110011111111100001001;
REG[8529] <= 32'b11110001111100110000000111111111;
REG[8530] <= 32'b11111100000100001111111100001101;
REG[8531] <= 32'b11110011000000010000000000000110;
REG[8532] <= 32'b00000001000101011110111111111111;
REG[8533] <= 32'b11111001000000111111011000001011;
REG[8534] <= 32'b11100111000001111111110000000101;
REG[8535] <= 32'b00000111000001010000110011101111;
REG[8536] <= 32'b11110011111101110001001000000001;
REG[8537] <= 32'b00010101111010111110100011101111;
REG[8538] <= 32'b00001010000001100001000011101101;
REG[8539] <= 32'b11110001111110111111101111111111;
REG[8540] <= 32'b00000100111101001111101111110011;
REG[8541] <= 32'b11111110111011101110110000001001;
REG[8542] <= 32'b00000101111101011111011011101110;
REG[8543] <= 32'b11110001111111001111000011110111;
REG[8544] <= 32'b11111010111101111111000011110100;
REG[8545] <= 32'b11111001000001111110111111110100;
REG[8546] <= 32'b11111010111011111111111000001011;
REG[8547] <= 32'b11110110111110101111000011110110;
REG[8548] <= 32'b11111110000010100000000100000000;
REG[8549] <= 32'b00000100111101001111100100000100;
REG[8550] <= 32'b00001001000001100000100000000011;
REG[8551] <= 32'b11110111000000000000001011111111;
REG[8552] <= 32'b11111110111101101111010111111101;
REG[8553] <= 32'b00000000111111000000001100000100;
REG[8554] <= 32'b00000101111110110000001111110011;
REG[8555] <= 32'b11111111001001010001000111110100;
REG[8556] <= 32'b00001010111111101111111111110101;
REG[8557] <= 32'b11111111111111000000011100000010;
REG[8558] <= 32'b11111111111110101111111000000000;
REG[8559] <= 32'b00000001111100001111110011110101;
REG[8560] <= 32'b11110110000001110000000011110011;
REG[8561] <= 32'b11111101111110101111101011111010;
REG[8562] <= 32'b11111000111111000000010000000110;
REG[8563] <= 32'b00000111000000101111010111111111;
REG[8564] <= 32'b00000000111111100000011111111000;
REG[8565] <= 32'b11101100000001001111011000000010;
REG[8566] <= 32'b00001011111111101111101011111110;
REG[8567] <= 32'b11111110000000001111011011111000;
REG[8568] <= 32'b11111110000010100000001000000110;
REG[8569] <= 32'b11111000111100011111011100000001;
REG[8570] <= 32'b11111001000011011111111011111000;
REG[8571] <= 32'b11111110111111110000001100000001;
REG[8572] <= 32'b00000101111111101111111000000000;
REG[8573] <= 32'b11111001111110110001010100000101;
REG[8574] <= 32'b11110111111101001111011011110101;
REG[8575] <= 32'b00010010111111111111000111111010;
REG[8576] <= 32'b11101110111101101111100000001010;
REG[8577] <= 32'b11111010000000011111000011111100;
REG[8578] <= 32'b11111011000001111111011011111100;
REG[8579] <= 32'b11110000000000000000000111111101;
REG[8580] <= 32'b11110111111011110000100000000011;
REG[8581] <= 32'b11111110000010001111011111110011;
REG[8582] <= 32'b00010010111110011111111100010000;
REG[8583] <= 32'b00001110000000010000111111111101;
REG[8584] <= 32'b00000111000110010000001011110101;
REG[8585] <= 32'b00000101000001110000000111111111;
REG[8586] <= 32'b11111110111010111111010100010101;
REG[8587] <= 32'b00000110000000010000100100000001;
REG[8588] <= 32'b00000111000011011111110011110110;
REG[8589] <= 32'b00000100000001011111111111111010;
REG[8590] <= 32'b11111111111101111111100000001000;
REG[8591] <= 32'b11110001111101010001011000000000;
REG[8592] <= 32'b11110001000001100000001011111101;
REG[8593] <= 32'b00001011000001001110110011101110;
REG[8594] <= 32'b00000001000010010000010000000010;
REG[8595] <= 32'b11111010111101001111011000000110;
REG[8596] <= 32'b00000011000010001111111011111110;
REG[8597] <= 32'b11110100000011100001000100001101;
REG[8598] <= 32'b11110100000001000000011100000000;
REG[8599] <= 32'b11111110111101101111001000000100;
REG[8600] <= 32'b00001000111101101111101011101101;
REG[8601] <= 32'b11111111111110011111100100000000;
REG[8602] <= 32'b11110011111101001111010011111000;
REG[8603] <= 32'b11111101111110011111100100000101;
REG[8604] <= 32'b11110011000001000000010111111101;
REG[8605] <= 32'b11111010000001101110101111110101;
REG[8606] <= 32'b11111000111111011111100100000001;
REG[8607] <= 32'b11111110111111010000011100000100;
REG[8608] <= 32'b00000101111111111111100000000000;
REG[8609] <= 32'b00001001000001010000101111111111;
REG[8610] <= 32'b00000101111111010000100000010000;
REG[8611] <= 32'b00010010000001000000101111111101;
REG[8612] <= 32'b11111101000010110000110100001011;
REG[8613] <= 32'b00011110000011111111111100000100;
REG[8614] <= 32'b00001001000001000001010111111111;
REG[8615] <= 32'b11111010000011010001001000001101;
REG[8616] <= 32'b11110100111001011111000000000011;
REG[8617] <= 32'b00010011111100101111011111100010;
REG[8618] <= 32'b11100101111101000001111000000100;
REG[8619] <= 32'b11111101111011101111011011111100;
REG[8620] <= 32'b00010101000001011111000111110001;
REG[8621] <= 32'b00000010111101010000010100000100;
REG[8622] <= 32'b11111001111101011111101000000010;
REG[8623] <= 32'b11111001111111001111110111111111;
REG[8624] <= 32'b00000001000000001111000011110100;
REG[8625] <= 32'b11101011000000000000001011111111;
REG[8626] <= 32'b00010000000010011111110000010011;
REG[8627] <= 32'b11111111000010010010110100001001;
REG[8628] <= 32'b11111101111111000000011011111010;
REG[8629] <= 32'b00010100000000000000100000001011;
REG[8630] <= 32'b00000101000011110000010011111111;
REG[8631] <= 32'b00000001000000010000010100011011;
REG[8632] <= 32'b11111010111111001111111011111100;
REG[8633] <= 32'b00000001000100111110111011110011;
REG[8634] <= 32'b11111110111100111111010011110011;
REG[8635] <= 32'b00000000000010111111000111101110;
REG[8636] <= 32'b11110001111100101111111000000010;
REG[8637] <= 32'b11111100111110011111011111110011;
REG[8638] <= 32'b11111011000000110000000100000100;
REG[8639] <= 32'b11100101000011010000011011111101;
REG[8640] <= 32'b00000110000010101111001100000010;
REG[8641] <= 32'b00001011000010010000010111111001;
REG[8642] <= 32'b11110001000010000000011111111100;
REG[8643] <= 32'b11111101000010111111101011111011;
REG[8644] <= 32'b00000000111111000000001000010001;
REG[8645] <= 32'b11110110000000010000011011111101;
REG[8646] <= 32'b11110011111101101111100111110111;
REG[8647] <= 32'b11111100111110101111001011111010;
REG[8648] <= 32'b11110100000000011111111011111010;
REG[8649] <= 32'b00001100000110000000101100000001;
REG[8650] <= 32'b11111101111110001111101100001110;
REG[8651] <= 32'b00000000111110001111110111110101;
REG[8652] <= 32'b11111010111110110000000000001111;
REG[8653] <= 32'b00000101000100100000000000000101;
REG[8654] <= 32'b00000111111111010000001000001101;
REG[8655] <= 32'b11101011111011001111110000010100;
REG[8656] <= 32'b00000110000011101111111011110011;
REG[8657] <= 32'b11110011000001001111110100000000;
REG[8658] <= 32'b11111100111100001110110111111100;
REG[8659] <= 32'b11111011000001011111101011110011;
REG[8660] <= 32'b11110111000001010000100000000011;
REG[8661] <= 32'b00000010000000110000000100001101;
REG[8662] <= 32'b11111000111101001111110011111011;
REG[8663] <= 32'b11110000000010110000010111111000;
REG[8664] <= 32'b00001100000000111111100100000001;
REG[8665] <= 32'b00010010111111011110011111111111;
REG[8666] <= 32'b00001111000001000000010000000111;
REG[8667] <= 32'b11110011000010010000100011111000;
REG[8668] <= 32'b11110011000001011111101100001101;
REG[8669] <= 32'b00001111000000001111001100000110;
REG[8670] <= 32'b11100111111101010000110000010101;
REG[8671] <= 32'b00000100111101101111000100001011;
REG[8672] <= 32'b00110101000010001111101011111000;
REG[8673] <= 32'b11111110000100010001010100010000;
REG[8674] <= 32'b11101110111110010000001011111100;
REG[8675] <= 32'b11101010111111111111111111111001;
REG[8676] <= 32'b00000000000001111110101011111101;
REG[8677] <= 32'b00001011000010111111101111111110;
REG[8678] <= 32'b11101111000000010000001100001000;
REG[8679] <= 32'b00000000000011101111111111111011;
REG[8680] <= 32'b11111011111101010000110000100100;
REG[8681] <= 32'b00001001111101010000101111111100;
REG[8682] <= 32'b00000101000100110000110011111110;
REG[8683] <= 32'b00000000111111110000100011110011;
REG[8684] <= 32'b11111101000010000000000011111101;
REG[8685] <= 32'b00000110111110000000001011111001;
REG[8686] <= 32'b11111010111111000000001011110101;
REG[8687] <= 32'b00000100000010110000010100000001;
REG[8688] <= 32'b11111110111101111111001111110100;
REG[8689] <= 32'b11110101111101100000110000001011;
REG[8690] <= 32'b00000001111110110000010100001101;
REG[8691] <= 32'b00000001111110001111110000000011;
REG[8692] <= 32'b00001010000010111110111000001110;
REG[8693] <= 32'b00000011000000101111101000001100;
REG[8694] <= 32'b00001110000110100000101011111111;
REG[8695] <= 32'b00000101000011100000110000010110;
REG[8696] <= 32'b00000000111111101111011011111110;
REG[8697] <= 32'b00000010111110000000010111111101;
REG[8698] <= 32'b00000000000011110000010011111100;
REG[8699] <= 32'b00010111000010100000010000000000;
REG[8700] <= 32'b11101101111100110000110111111001;
REG[8701] <= 32'b00000101000011010000110000000101;
REG[8702] <= 32'b00000000111111100001010000001100;
REG[8703] <= 32'b11101101111100011111011000000001;
REG[8704] <= 32'b00010101000010011111000111101010;
REG[8705] <= 32'b00001001111110010000111011111000;
REG[8706] <= 32'b11110010111100000000001100000000;
REG[8707] <= 32'b11110110111101011111010011110110;
REG[8708] <= 32'b00000001111110100000000000000100;
REG[8709] <= 32'b11110100111101111111110011101110;
REG[8710] <= 32'b00000101000010100000001111111010;
REG[8711] <= 32'b11111110000000011111100100000110;
REG[8712] <= 32'b00000000111100111111100111111101;
REG[8713] <= 32'b11111101111111101110101011110001;
REG[8714] <= 32'b11111101000000101111111100000000;
REG[8715] <= 32'b00000001000010111111110111111011;
REG[8716] <= 32'b11111001000010000000100100001000;
REG[8717] <= 32'b11110110000001010000011000000100;
REG[8718] <= 32'b00010011000001111111000100000001;
REG[8719] <= 32'b00001110000001010000100000001101;
REG[8720] <= 32'b00001111111110001111011111111011;
REG[8721] <= 32'b11111111111101110001011100101111;
REG[8722] <= 32'b00100011000000010001011100011100;
REG[8723] <= 32'b00011101111101001111110011111110;
REG[8724] <= 32'b00000100000001110000000011110100;
REG[8725] <= 32'b11101000000000100000010011111001;
REG[8726] <= 32'b11110111000010001110111111111111;
REG[8727] <= 32'b11111011111100110000101011111111;
REG[8728] <= 32'b11101111000001110000111111110000;
REG[8729] <= 32'b00001001000001100000000111101111;
REG[8730] <= 32'b00010100111100101111100000010010;
REG[8731] <= 32'b00100010000000110000001000000010;
REG[8732] <= 32'b00001010111100100000011111110011;
REG[8733] <= 32'b00001101111111111111101100000101;
REG[8734] <= 32'b00001010000010110000000111110110;
REG[8735] <= 32'b11111001111111100000010111111010;
REG[8736] <= 32'b11111111111101111111111000000110;
REG[8737] <= 32'b00001101000000111110101100000010;
REG[8738] <= 32'b11110101111111111111100011101011;
REG[8739] <= 32'b11111011000001011111101011111010;
REG[8740] <= 32'b00001001000001000000011100000100;
REG[8741] <= 32'b11111000000001000000011000000101;
REG[8742] <= 32'b00010010000100010000001011111110;
REG[8743] <= 32'b00000000000001110001111100100110;
REG[8744] <= 32'b00001100111111110000001100000111;
REG[8745] <= 32'b11110101000011111111011000000000;
REG[8746] <= 32'b11111010111110111110111000000000;
REG[8747] <= 32'b00001101000011010000111100001110;
REG[8748] <= 32'b00010101001000000000001000001011;
REG[8749] <= 32'b00000011000001101110000100010010;
REG[8750] <= 32'b11111110000001010000011000000111;
REG[8751] <= 32'b00001001111101111111001011111010;
REG[8752] <= 32'b11111001111110011111111011101111;
REG[8753] <= 32'b11110001111101001111011100000000;
REG[8754] <= 32'b00001000111101011111010011111011;
REG[8755] <= 32'b11111000111111011111011011111011;
REG[8756] <= 32'b00010011000000111111100111111000;
REG[8757] <= 32'b11111101000001010000001111111111;
REG[8758] <= 32'b11110111000001001111011111110011;
REG[8759] <= 32'b11110001000101000000001100000110;
REG[8760] <= 32'b00010100111111011111010111111100;
REG[8761] <= 32'b11110011000000000000111111111111;
REG[8762] <= 32'b11110011111010011110001011110100;
REG[8763] <= 32'b00011110000111111111110011110000;
REG[8764] <= 32'b11011101111110011110101111111000;
REG[8765] <= 32'b11110001111111101111101100000101;
REG[8766] <= 32'b11111101000010101111101100001100;
REG[8767] <= 32'b00010010000100101110010000010011;
REG[8768] <= 32'b00000000111111110000010000001000;
REG[8769] <= 32'b11111000111111101111111100000011;
REG[8770] <= 32'b00000001000000111111111111111110;
REG[8771] <= 32'b00000010000000000000000111110100;
REG[8772] <= 32'b11111011111110111111111100001010;
REG[8773] <= 32'b11111101111111011111001111111001;
REG[8774] <= 32'b11111101111111101111111100000000;
REG[8775] <= 32'b11111100111110101110111000000000;
REG[8776] <= 32'b11111100111101100001010111111101;
REG[8777] <= 32'b11110110111111111111111111111110;
REG[8778] <= 32'b11111010000100100001011111110110;
REG[8779] <= 32'b00000110000001000001001100001011;
REG[8780] <= 32'b11111110111111010001001000001010;
REG[8781] <= 32'b00011000000010111111000111110100;
REG[8782] <= 32'b00001000000000101111011011111001;
REG[8783] <= 32'b11110100111111010000000100000101;
REG[8784] <= 32'b00010111000100110000100111111011;
REG[8785] <= 32'b00000111000001100000010111110101;
REG[8786] <= 32'b11100001000001000000101100000111;
REG[8787] <= 32'b00000100111111011111111111111111;
REG[8788] <= 32'b00000100000000010000011000000101;
REG[8789] <= 32'b00000001111110010000011100001010;
REG[8790] <= 32'b00001111111111100000001011111101;
REG[8791] <= 32'b00000111000011110000110000000000;
REG[8792] <= 32'b00001100111111001111101011111000;
REG[8793] <= 32'b00000101000000000000111100100100;
REG[8794] <= 32'b00010011111111011111111011111101;
REG[8795] <= 32'b11111000000100010000101000000010;
REG[8796] <= 32'b00001001111110110000010011110110;
REG[8797] <= 32'b11111100111110000000011100000101;
REG[8798] <= 32'b11111110111101111111101011110001;
REG[8799] <= 32'b11111010111110100000010011111010;
REG[8800] <= 32'b11110010111010110000101100100101;
REG[8801] <= 32'b00000011000010000001001011111101;
REG[8802] <= 32'b11111110111111100001110000000001;
REG[8803] <= 32'b00100001000010000000000100000000;
REG[8804] <= 32'b00001100000001110001011100000011;
REG[8805] <= 32'b11101010111111010000000000001000;
REG[8806] <= 32'b11111100111111000000001100000100;
REG[8807] <= 32'b11110010000001110000011111110111;
REG[8808] <= 32'b11111001111111001111011100001100;
REG[8809] <= 32'b00001000111101011111110011110111;
REG[8810] <= 32'b11101001000001110001010000010110;
REG[8811] <= 32'b00010110000001111110000100000100;
REG[8812] <= 32'b00001101000000100000101000001111;
REG[8813] <= 32'b11101011111111110000110000000100;
REG[8814] <= 32'b00000010111111110000010111101101;
REG[8815] <= 32'b11111110000000011111001111101111;
REG[8816] <= 32'b11111000000011010000000011111000;
REG[8817] <= 32'b00000011000000100000011000001010;
REG[8818] <= 32'b11111011111101111111100111111110;
REG[8819] <= 32'b11111111000001111111111111111111;
REG[8820] <= 32'b11110100000011010000000011110101;
REG[8821] <= 32'b11111100111101110000011011111010;
REG[8822] <= 32'b11111000111111111111111100000101;
REG[8823] <= 32'b11111101111101001111110111111110;
REG[8824] <= 32'b11111111111111011111011011101110;
REG[8825] <= 32'b11110100111101001111100011110110;
REG[8826] <= 32'b11111100111101001111011111111000;
REG[8827] <= 32'b11111101111111001111101011111111;
REG[8828] <= 32'b00010011111110100000101011110111;
REG[8829] <= 32'b11110110111100011111101111111000;
REG[8830] <= 32'b00000001111101101110010111101110;
REG[8831] <= 32'b11110100000010100000101111111010;
REG[8832] <= 32'b00000010111111000000001000000011;
REG[8833] <= 32'b00000100000000010000000000000010;
REG[8834] <= 32'b11111100111110000000001000000110;
REG[8835] <= 32'b11111001000000001111110011110111;
REG[8836] <= 32'b00000001000000010000001100000001;
REG[8837] <= 32'b00000000111111011111100000001001;
REG[8838] <= 32'b00000010000001110000000000000001;
REG[8839] <= 32'b11110111111111010001010100000100;
REG[8840] <= 32'b00000100111110101111001011101111;
REG[8841] <= 32'b11111100111101101111101011011001;
REG[8842] <= 32'b11100110000001110000010000000111;
REG[8843] <= 32'b00010011110101101111010100100100;
REG[8844] <= 32'b00000000000001000000011011101111;
REG[8845] <= 32'b11101100111111110000100100000101;
REG[8846] <= 32'b00001111000011010000111011110001;
REG[8847] <= 32'b00010001000000010000110111111001;
REG[8848] <= 32'b00000011000010110000110000000011;
REG[8849] <= 32'b00000001000010000000001000000100;
REG[8850] <= 32'b11111101111111001111011100000101;
REG[8851] <= 32'b00000101111100110000110000001101;
REG[8852] <= 32'b00000100111101001111100011110110;
REG[8853] <= 32'b00001010000100110000000011111001;
REG[8854] <= 32'b00000000111101111111110011110000;
REG[8855] <= 32'b11110110111100101111000111111010;
REG[8856] <= 32'b00001001111011101111011011111010;
REG[8857] <= 32'b11111111111101011111101011110000;
REG[8858] <= 32'b11110011111101010000001111111010;
REG[8859] <= 32'b00000101000001001111101011111101;
REG[8860] <= 32'b00000011111110000000010000001100;
REG[8861] <= 32'b00000100111111001111101111101111;
REG[8862] <= 32'b00000111000000111111110000000011;
REG[8863] <= 32'b00001000000000010000000011111111;
REG[8864] <= 32'b00000000000000010000010000000100;
REG[8865] <= 32'b00000011000010000000010011110101;
REG[8866] <= 32'b11111011000000110000011100001000;
REG[8867] <= 32'b00001000111110011111110000000101;
REG[8868] <= 32'b11111011111110110000001011111001;
REG[8869] <= 32'b11110100111111111111110011110111;
REG[8870] <= 32'b00001110000000111111100000001010;
REG[8871] <= 32'b00000000111110010000011011111011;
REG[8872] <= 32'b00000001000011011111100111101110;
REG[8873] <= 32'b00001011111100010000100000000111;
REG[8874] <= 32'b11110010111110010001011011111001;
REG[8875] <= 32'b11111011111101000000101000001100;
REG[8876] <= 32'b00011100000000001111111011110101;
REG[8877] <= 32'b00000001000001010000001000001110;
REG[8878] <= 32'b00000100000001010000101011111111;
REG[8879] <= 32'b11111001000011111111110011110010;
REG[8880] <= 32'b00000110111110111111100000000100;
REG[8881] <= 32'b11111011111101010000010011111011;
REG[8882] <= 32'b11110110111110110000011000010000;
REG[8883] <= 32'b00010000000000101111010011111010;
REG[8884] <= 32'b11111000111100110000101011111010;
REG[8885] <= 32'b11110101111110101111000111101110;
REG[8886] <= 32'b11111001000001000000100011111011;
REG[8887] <= 32'b00000011000010110000100000010101;
REG[8888] <= 32'b00100011111010111111011000001001;
REG[8889] <= 32'b11111001111110001111110111110111;
REG[8890] <= 32'b00001000000011111111011111111111;
REG[8891] <= 32'b11101000111110000000011111111011;
REG[8892] <= 32'b11111111000001011110110000000000;
REG[8893] <= 32'b00000111000001111111011011110110;
REG[8894] <= 32'b11110010111110100000011100001001;
REG[8895] <= 32'b00001110000000000000010011110101;
REG[8896] <= 32'b11111001111111010000101111111010;
REG[8897] <= 32'b11111010111001101110110011110010;
REG[8898] <= 32'b00001011000000010000010111110110;
REG[8899] <= 32'b11110001111110011111111011111111;
REG[8900] <= 32'b00000010000001010000000111111000;
REG[8901] <= 32'b00000010000001111111011111111100;
REG[8902] <= 32'b11111001111101101111111111111000;
REG[8903] <= 32'b11110101000001000000000011111010;
REG[8904] <= 32'b00000010111110111111111000000011;
REG[8905] <= 32'b00010001000010110001100000001001;
REG[8906] <= 32'b11111110111110100001000100001011;
REG[8907] <= 32'b00001111000000011111100000000100;
REG[8908] <= 32'b00001110000011110000000011111001;
REG[8909] <= 32'b11101011111100101111110100000011;
REG[8910] <= 32'b00000010111111001111110000000111;
REG[8911] <= 32'b11111110111100001111101111110101;
REG[8912] <= 32'b11110011000001110000000011111000;
REG[8913] <= 32'b11110000111100101111110011111010;
REG[8914] <= 32'b11111001111110101111101011110111;
REG[8915] <= 32'b00000100000010001111011011110101;
REG[8916] <= 32'b00000001000001110001011000000011;
REG[8917] <= 32'b00000101111111011111100011111101;
REG[8918] <= 32'b00001000000011100001001000010101;
REG[8919] <= 32'b00001000000000000000100111111101;
REG[8920] <= 32'b11111101000011001111101111111100;
REG[8921] <= 32'b00001010111101101111011100000111;
REG[8922] <= 32'b11111011111111011111110000000010;
REG[8923] <= 32'b00100111000101111111100100000011;
REG[8924] <= 32'b11111111000100010010011111111110;
REG[8925] <= 32'b11110000000000110000001100010101;
REG[8926] <= 32'b00011000111011011111111111111010;
REG[8927] <= 32'b11111011000000110000101111111111;
REG[8928] <= 32'b11111001111110011111010111111011;
REG[8929] <= 32'b11111100111100101111101111111101;
REG[8930] <= 32'b11111110111101001110111111110111;
REG[8931] <= 32'b00000010111111001111100000100000;
REG[8932] <= 32'b00001100000010011111111011111001;
REG[8933] <= 32'b11111000000111000000011111111001;
REG[8934] <= 32'b11110111111111111111101100001101;
REG[8935] <= 32'b00000101111100010000001000010010;
REG[8936] <= 32'b00000001000101010000001100000000;
REG[8937] <= 32'b00001111000100101111110000010000;
REG[8938] <= 32'b00001010000001111111110011111110;
REG[8939] <= 32'b11110010111111000000010000000100;
REG[8940] <= 32'b11111110111110010000011100000011;
REG[8941] <= 32'b11111110000010111111100111110110;
REG[8942] <= 32'b11111111000010011111110111110110;
REG[8943] <= 32'b00000000111111110000100100000011;
REG[8944] <= 32'b00000110000000111111110000000101;
REG[8945] <= 32'b11111100111110111111010011111100;
REG[8946] <= 32'b11110110000001000000011000001111;
REG[8947] <= 32'b00000110000001011111001111110110;
REG[8948] <= 32'b11111101111111001111100100010011;
REG[8949] <= 32'b11111100111110101111111111101100;
REG[8950] <= 32'b00000001001110111111011111110001;
REG[8951] <= 32'b00000000111100111111100000001110;
REG[8952] <= 32'b11111010111101111111011111110001;
REG[8953] <= 32'b11111001000010010000001000000000;
REG[8954] <= 32'b00000001111111011111101111111100;
REG[8955] <= 32'b00000011111110010000011100000011;
REG[8956] <= 32'b11111110000000011111111111111110;
REG[8957] <= 32'b00000001000010010000001000000110;
REG[8958] <= 32'b11111110000001111111111111111110;
REG[8959] <= 32'b00000111111101000000000000010100;
REG[8960] <= 32'b00001100111010100001001111110100;
REG[8961] <= 32'b11111011000000001111111111111001;
REG[8962] <= 32'b00010010111110100000110100010001;
REG[8963] <= 32'b11111000000000110000001100010011;
REG[8964] <= 32'b00100011000111101111100011101010;
REG[8965] <= 32'b11111101111100110000010011110111;
REG[8966] <= 32'b11110000111110010000110111111110;
REG[8967] <= 32'b11111100111111100000010011111100;
REG[8968] <= 32'b00000010000000100000001000000101;
REG[8969] <= 32'b00001010111100111111001111110101;
REG[8970] <= 32'b00000111000001010000101011111010;
REG[8971] <= 32'b11101110111110000000110000001011;
REG[8972] <= 32'b00001011111110110000000100000010;
REG[8973] <= 32'b00001010000011011111110111111000;
REG[8974] <= 32'b11110111111101110000001011111001;
REG[8975] <= 32'b11111011111100001111011011110111;


	end
	else if(i_wr_en) begin
		REG[i_wr_addr] <= i_wr_data; // Write behavior
	end
end

endmodule